/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
****************************************************************************
*
* Module    : wav_mcuintf_csr_defs.vh
* Date      : 2021-01-14
* Desciption: Autogenerated CSR block.
*
* $Id: wav_mcuintf_csr_defs.vh,v 1.6 2021/01/15 11:30:08 schilukuri Exp $
*
****************************************************************************/

// Word Address 0x00000000 : WAV_MCUINTF_HOST2MCU_MSG_DATA (RW)
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_DATA_FIELD 31:0
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_DATA_FIELD_WIDTH 32
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_RANGE 31:0
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_WIDTH 32
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_ADR 32'h00000000
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_POR 32'h00000000
`define WAV_MCUINTF_HOST2MCU_MSG_DATA_MSK 32'hFFFFFFFF

// Word Address 0x00000004 : WAV_MCUINTF_HOST2MCU_MSG_ID (RW)
`define WAV_MCUINTF_HOST2MCU_MSG_ID_ID_FIELD 31:0
`define WAV_MCUINTF_HOST2MCU_MSG_ID_ID_FIELD_WIDTH 32
`define WAV_MCUINTF_HOST2MCU_MSG_ID_RANGE 31:0
`define WAV_MCUINTF_HOST2MCU_MSG_ID_WIDTH 32
`define WAV_MCUINTF_HOST2MCU_MSG_ID_ADR 32'h00000004
`define WAV_MCUINTF_HOST2MCU_MSG_ID_POR 32'h00000000
`define WAV_MCUINTF_HOST2MCU_MSG_ID_MSK 32'hFFFFFFFF

// Word Address 0x00000008 : WAV_MCUINTF_HOST2MCU_MSG_REQ (W1T)
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_REQ_FIELD 0
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_REQ_FIELD_WIDTH 1
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_RANGE 0:0
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_WIDTH 1
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_ADR 32'h00000008
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_POR 32'h00000000
`define WAV_MCUINTF_HOST2MCU_MSG_REQ_MSK 32'h00000001

// Word Address 0x0000000C : WAV_MCUINTF_HOST2MCU_MSG_ACK (W1T)
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_ACK_FIELD 0
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_ACK_FIELD_WIDTH 1
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_RANGE 0:0
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_WIDTH 1
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_ADR 32'h0000000C
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_POR 32'h00000000
`define WAV_MCUINTF_HOST2MCU_MSG_ACK_MSK 32'h00000001

// Word Address 0x00000010 : WAV_MCUINTF_MCU2HOST_MSG_DATA (RW)
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_DATA_FIELD 31:0
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_DATA_FIELD_WIDTH 32
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_RANGE 31:0
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_WIDTH 32
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_ADR 32'h00000010
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_POR 32'h00000000
`define WAV_MCUINTF_MCU2HOST_MSG_DATA_MSK 32'hFFFFFFFF

// Word Address 0x00000014 : WAV_MCUINTF_MCU2HOST_MSG_ID (RW)
`define WAV_MCUINTF_MCU2HOST_MSG_ID_ID_FIELD 31:0
`define WAV_MCUINTF_MCU2HOST_MSG_ID_ID_FIELD_WIDTH 32
`define WAV_MCUINTF_MCU2HOST_MSG_ID_RANGE 31:0
`define WAV_MCUINTF_MCU2HOST_MSG_ID_WIDTH 32
`define WAV_MCUINTF_MCU2HOST_MSG_ID_ADR 32'h00000014
`define WAV_MCUINTF_MCU2HOST_MSG_ID_POR 32'h00000000
`define WAV_MCUINTF_MCU2HOST_MSG_ID_MSK 32'hFFFFFFFF

// Word Address 0x00000018 : WAV_MCUINTF_MCU2HOST_MSG_REQ (W1T)
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_REQ_FIELD 0
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_REQ_FIELD_WIDTH 1
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_RANGE 0:0
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_WIDTH 1
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_ADR 32'h00000018
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_POR 32'h00000000
`define WAV_MCUINTF_MCU2HOST_MSG_REQ_MSK 32'h00000001

// Word Address 0x0000001C : WAV_MCUINTF_MCU2HOST_MSG_ACK (W1T)
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_ACK_FIELD 0
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_ACK_FIELD_WIDTH 1
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_RANGE 0:0
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_WIDTH 1
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_ADR 32'h0000001C
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_POR 32'h00000000
`define WAV_MCUINTF_MCU2HOST_MSG_ACK_MSK 32'h00000001
