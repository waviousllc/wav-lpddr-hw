/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
****************************************************************************
*
* Module    : ddr_fsw_csr_defs.vh
* Date      : 2021-04-22
* Desciption: Autogenerated CSR block.
*
* $Id: ddr_fsw_csr_defs.vh,v 1.35 2021/04/23 22:16:09 mclovis Exp $
*
****************************************************************************/

// Word Address 0x00000000 : DDR_FSW_CTRL_CFG (RW)
`define DDR_FSW_CTRL_CFG_MSR_OVR_FIELD 6
`define DDR_FSW_CTRL_CFG_MSR_OVR_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_MSR_OVR_VAL_FIELD 7
`define DDR_FSW_CTRL_CFG_MSR_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_MSR_TOGGLE_EN_FIELD 5
`define DDR_FSW_CTRL_CFG_MSR_TOGGLE_EN_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_POST_GFMSEL_WAIT_FIELD 19:16
`define DDR_FSW_CTRL_CFG_POST_GFMSEL_WAIT_FIELD_WIDTH 4
`define DDR_FSW_CTRL_CFG_PREP_DONE_FIELD 8
`define DDR_FSW_CTRL_CFG_PREP_DONE_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_PSTWORK_DONE_FIELD 9
`define DDR_FSW_CTRL_CFG_PSTWORK_DONE_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_PSTWORK_DONE_OVR_FIELD 10
`define DDR_FSW_CTRL_CFG_PSTWORK_DONE_OVR_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_SWITCH_DONE_OVR_FIELD 11
`define DDR_FSW_CTRL_CFG_SWITCH_DONE_OVR_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_SWITCH_DONE_STICKY_CLR_FIELD 12
`define DDR_FSW_CTRL_CFG_SWITCH_DONE_STICKY_CLR_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_VCO_SEL_OVR_FIELD 0
`define DDR_FSW_CTRL_CFG_VCO_SEL_OVR_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_VCO_SEL_OVR_VAL_FIELD 2:1
`define DDR_FSW_CTRL_CFG_VCO_SEL_OVR_VAL_FIELD_WIDTH 2
`define DDR_FSW_CTRL_CFG_VCO_TOGGLE_EN_FIELD 4
`define DDR_FSW_CTRL_CFG_VCO_TOGGLE_EN_FIELD_WIDTH 1
`define DDR_FSW_CTRL_CFG_RANGE 19:0
`define DDR_FSW_CTRL_CFG_WIDTH 20
`define DDR_FSW_CTRL_CFG_ADR 32'h00000000
`define DDR_FSW_CTRL_CFG_POR 32'h00040C31
`define DDR_FSW_CTRL_CFG_MSK 32'h000F1FF7

// Word Address 0x00000004 : DDR_FSW_CTRL_STA (R)
`define DDR_FSW_CTRL_STA_CMN_MSR_FIELD 3
`define DDR_FSW_CTRL_STA_CMN_MSR_FIELD_WIDTH 1
`define DDR_FSW_CTRL_STA_CORE_READY_FIELD 4
`define DDR_FSW_CTRL_STA_CORE_READY_FIELD_WIDTH 1
`define DDR_FSW_CTRL_STA_SWITCH_DONE_FIELD 2
`define DDR_FSW_CTRL_STA_SWITCH_DONE_FIELD_WIDTH 1
`define DDR_FSW_CTRL_STA_VCO_SEL_FIELD 1:0
`define DDR_FSW_CTRL_STA_VCO_SEL_FIELD_WIDTH 2
`define DDR_FSW_CTRL_STA_RANGE 4:0
`define DDR_FSW_CTRL_STA_WIDTH 5
`define DDR_FSW_CTRL_STA_ADR 32'h00000004
`define DDR_FSW_CTRL_STA_POR 32'h00000000
`define DDR_FSW_CTRL_STA_MSK 32'h0000001F

// Word Address 0x00000008 : DDR_FSW_DEBUG_CFG (RW)
`define DDR_FSW_DEBUG_CFG_DEBUG_BUS_SEL_FIELD 3:0
`define DDR_FSW_DEBUG_CFG_DEBUG_BUS_SEL_FIELD_WIDTH 4
`define DDR_FSW_DEBUG_CFG_RANGE 3:0
`define DDR_FSW_DEBUG_CFG_WIDTH 4
`define DDR_FSW_DEBUG_CFG_ADR 32'h00000008
`define DDR_FSW_DEBUG_CFG_POR 32'h00000000
`define DDR_FSW_DEBUG_CFG_MSK 32'h0000000F

// Word Address 0x0000002C : DDR_FSW_CSP_0_CFG (RW)
`define DDR_FSW_CSP_0_CFG_PRECLKDIS_WAIT_FIELD 3:0
`define DDR_FSW_CSP_0_CFG_PRECLKDIS_WAIT_FIELD_WIDTH 4
`define DDR_FSW_CSP_0_CFG_PRERST_WAIT_FIELD 7:4
`define DDR_FSW_CSP_0_CFG_PRERST_WAIT_FIELD_WIDTH 4
`define DDR_FSW_CSP_0_CFG_PSTCLKEN_WAIT_FIELD 19:16
`define DDR_FSW_CSP_0_CFG_PSTCLKEN_WAIT_FIELD_WIDTH 4
`define DDR_FSW_CSP_0_CFG_PSTPIEN_WAIT_FIELD 23:20
`define DDR_FSW_CSP_0_CFG_PSTPIEN_WAIT_FIELD_WIDTH 4
`define DDR_FSW_CSP_0_CFG_PSTRST_WAIT_FIELD 15:12
`define DDR_FSW_CSP_0_CFG_PSTRST_WAIT_FIELD_WIDTH 4
`define DDR_FSW_CSP_0_CFG_RST_PULSE_WIDTH_FIELD 11:8
`define DDR_FSW_CSP_0_CFG_RST_PULSE_WIDTH_FIELD_WIDTH 4
`define DDR_FSW_CSP_0_CFG_RANGE 23:0
`define DDR_FSW_CSP_0_CFG_WIDTH 24
`define DDR_FSW_CSP_0_CFG_ADR 32'h0000002C
`define DDR_FSW_CSP_0_CFG_POR 32'h00333333
`define DDR_FSW_CSP_0_CFG_MSK 32'h00FFFFFF

// Word Address 0x00000030 : DDR_FSW_CSP_1_CFG (RW)
`define DDR_FSW_CSP_1_CFG_CGC_EN_OVR_FIELD 2
`define DDR_FSW_CSP_1_CFG_CGC_EN_OVR_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_CGC_EN_OVR_VAL_FIELD 5
`define DDR_FSW_CSP_1_CFG_CGC_EN_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_CLK_DISABLE_OVR_VAL_FIELD 8
`define DDR_FSW_CSP_1_CFG_CLK_DISABLE_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_DIV_RST_OVR_VAL_FIELD 7
`define DDR_FSW_CSP_1_CFG_DIV_RST_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_PI_DISABLE_OVR_VAL_FIELD 6
`define DDR_FSW_CSP_1_CFG_PI_DISABLE_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_REQ_COMPLETE_OVR_FIELD 1
`define DDR_FSW_CSP_1_CFG_REQ_COMPLETE_OVR_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_REQ_COMPLETE_OVR_VAL_FIELD 4
`define DDR_FSW_CSP_1_CFG_REQ_COMPLETE_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_REQ_COMPLETE_STA_CLR_FIELD 9
`define DDR_FSW_CSP_1_CFG_REQ_COMPLETE_STA_CLR_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_REQ_OVR_FIELD 0
`define DDR_FSW_CSP_1_CFG_REQ_OVR_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_REQ_OVR_VAL_FIELD 3
`define DDR_FSW_CSP_1_CFG_REQ_OVR_VAL_FIELD_WIDTH 1
`define DDR_FSW_CSP_1_CFG_RANGE 9:0
`define DDR_FSW_CSP_1_CFG_WIDTH 10
`define DDR_FSW_CSP_1_CFG_ADR 32'h00000030
`define DDR_FSW_CSP_1_CFG_POR 32'h00000100
`define DDR_FSW_CSP_1_CFG_MSK 32'h000003FF

// Word Address 0x00000034 : DDR_FSW_CSP_STA (R)
`define DDR_FSW_CSP_STA_REQ_COMPLETE_FIELD 0
`define DDR_FSW_CSP_STA_REQ_COMPLETE_FIELD_WIDTH 1
`define DDR_FSW_CSP_STA_RANGE 0:0
`define DDR_FSW_CSP_STA_WIDTH 1
`define DDR_FSW_CSP_STA_ADR 32'h00000034
`define DDR_FSW_CSP_STA_POR 32'h00000000
`define DDR_FSW_CSP_STA_MSK 32'h00000001
