/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
****************************************************************************
*
* Module    : ddr_cmn_csr_defs.vh
* Date      : 2021-04-22
* Desciption: Autogenerated CSR block.
*
* $Id: ddr_cmn_csr_defs.vh,v 1.149 2021/04/23 22:16:09 mclovis Exp $
*
****************************************************************************/

// Word Address 0x00000008 : DDR_CMN_VREF_M0_CFG (RW)
`define DDR_CMN_VREF_M0_CFG_CTRL_FIELD 7:0
`define DDR_CMN_VREF_M0_CFG_CTRL_FIELD_WIDTH 8
`define DDR_CMN_VREF_M0_CFG_EN_FIELD 9
`define DDR_CMN_VREF_M0_CFG_EN_FIELD_WIDTH 1
`define DDR_CMN_VREF_M0_CFG_HIZ_FIELD 10
`define DDR_CMN_VREF_M0_CFG_HIZ_FIELD_WIDTH 1
`define DDR_CMN_VREF_M0_CFG_PWR_FIELD 12:11
`define DDR_CMN_VREF_M0_CFG_PWR_FIELD_WIDTH 2
`define DDR_CMN_VREF_M0_CFG_RANGE 12:0
`define DDR_CMN_VREF_M0_CFG_WIDTH 13
`define DDR_CMN_VREF_M0_CFG_ADR 32'h00000008
`define DDR_CMN_VREF_M0_CFG_POR 32'h00000000
`define DDR_CMN_VREF_M0_CFG_MSK 32'h00001EFF

// Word Address 0x0000000C : DDR_CMN_VREF_M1_CFG (RW)
`define DDR_CMN_VREF_M1_CFG_CTRL_FIELD 7:0
`define DDR_CMN_VREF_M1_CFG_CTRL_FIELD_WIDTH 8
`define DDR_CMN_VREF_M1_CFG_EN_FIELD 9
`define DDR_CMN_VREF_M1_CFG_EN_FIELD_WIDTH 1
`define DDR_CMN_VREF_M1_CFG_HIZ_FIELD 10
`define DDR_CMN_VREF_M1_CFG_HIZ_FIELD_WIDTH 1
`define DDR_CMN_VREF_M1_CFG_PWR_FIELD 12:11
`define DDR_CMN_VREF_M1_CFG_PWR_FIELD_WIDTH 2
`define DDR_CMN_VREF_M1_CFG_RANGE 12:0
`define DDR_CMN_VREF_M1_CFG_WIDTH 13
`define DDR_CMN_VREF_M1_CFG_ADR 32'h0000000C
`define DDR_CMN_VREF_M1_CFG_POR 32'h00000000
`define DDR_CMN_VREF_M1_CFG_MSK 32'h00001EFF

// Word Address 0x00000010 : DDR_CMN_ZQCAL_CFG (RW)
`define DDR_CMN_ZQCAL_CFG_CAL_EN_FIELD 5
`define DDR_CMN_ZQCAL_CFG_CAL_EN_FIELD_WIDTH 1
`define DDR_CMN_ZQCAL_CFG_NCAL_FIELD 4:0
`define DDR_CMN_ZQCAL_CFG_NCAL_FIELD_WIDTH 5
`define DDR_CMN_ZQCAL_CFG_PCAL_FIELD 13:8
`define DDR_CMN_ZQCAL_CFG_PCAL_FIELD_WIDTH 6
`define DDR_CMN_ZQCAL_CFG_PD_SEL_FIELD 6
`define DDR_CMN_ZQCAL_CFG_PD_SEL_FIELD_WIDTH 1
`define DDR_CMN_ZQCAL_CFG_VOL_0P6_SEL_FIELD 7
`define DDR_CMN_ZQCAL_CFG_VOL_0P6_SEL_FIELD_WIDTH 1
`define DDR_CMN_ZQCAL_CFG_RANGE 13:0
`define DDR_CMN_ZQCAL_CFG_WIDTH 14
`define DDR_CMN_ZQCAL_CFG_ADR 32'h00000010
`define DDR_CMN_ZQCAL_CFG_POR 32'h00000000
`define DDR_CMN_ZQCAL_CFG_MSK 32'h00003FFF

// Word Address 0x00000014 : DDR_CMN_ZQCAL_STA (R)
`define DDR_CMN_ZQCAL_STA_COMP_FIELD 0
`define DDR_CMN_ZQCAL_STA_COMP_FIELD_WIDTH 1
`define DDR_CMN_ZQCAL_STA_RANGE 0:0
`define DDR_CMN_ZQCAL_STA_WIDTH 1
`define DDR_CMN_ZQCAL_STA_ADR 32'h00000014
`define DDR_CMN_ZQCAL_STA_POR 32'h00000000
`define DDR_CMN_ZQCAL_STA_MSK 32'h00000001

// Word Address 0x00000018 : DDR_CMN_IBIAS_CFG (RW)
`define DDR_CMN_IBIAS_CFG_EN_FIELD 0
`define DDR_CMN_IBIAS_CFG_EN_FIELD_WIDTH 1
`define DDR_CMN_IBIAS_CFG_RANGE 0:0
`define DDR_CMN_IBIAS_CFG_WIDTH 1
`define DDR_CMN_IBIAS_CFG_ADR 32'h00000018
`define DDR_CMN_IBIAS_CFG_POR 32'h00000000
`define DDR_CMN_IBIAS_CFG_MSK 32'h00000001

// Word Address 0x0000001C : DDR_CMN_TEST_CFG (RW)
`define DDR_CMN_TEST_CFG_ATB_MODE_FIELD 1:0
`define DDR_CMN_TEST_CFG_ATB_MODE_FIELD_WIDTH 2
`define DDR_CMN_TEST_CFG_ATST_SEL_FIELD 5:2
`define DDR_CMN_TEST_CFG_ATST_SEL_FIELD_WIDTH 4
`define DDR_CMN_TEST_CFG_DTST_DIV_EN_FIELD 17
`define DDR_CMN_TEST_CFG_DTST_DIV_EN_FIELD_WIDTH 1
`define DDR_CMN_TEST_CFG_DTST_DRVR_IMPD_FIELD 10:8
`define DDR_CMN_TEST_CFG_DTST_DRVR_IMPD_FIELD_WIDTH 3
`define DDR_CMN_TEST_CFG_DTST_EXT_SEL_FIELD 16:12
`define DDR_CMN_TEST_CFG_DTST_EXT_SEL_FIELD_WIDTH 5
`define DDR_CMN_TEST_CFG_RANGE 17:0
`define DDR_CMN_TEST_CFG_WIDTH 18
`define DDR_CMN_TEST_CFG_ADR 32'h0000001C
`define DDR_CMN_TEST_CFG_POR 32'h00000000
`define DDR_CMN_TEST_CFG_MSK 32'h0003F73F

// Word Address 0x00000020 : DDR_CMN_LDO_M0_CFG (RW)
`define DDR_CMN_LDO_M0_CFG_ATST_SEL_FIELD 12:10
`define DDR_CMN_LDO_M0_CFG_ATST_SEL_FIELD_WIDTH 3
`define DDR_CMN_LDO_M0_CFG_EN_FIELD 8
`define DDR_CMN_LDO_M0_CFG_EN_FIELD_WIDTH 1
`define DDR_CMN_LDO_M0_CFG_HIZ_FIELD 13
`define DDR_CMN_LDO_M0_CFG_HIZ_FIELD_WIDTH 1
`define DDR_CMN_LDO_M0_CFG_TRAN_ENH_EN_FIELD 9
`define DDR_CMN_LDO_M0_CFG_TRAN_ENH_EN_FIELD_WIDTH 1
`define DDR_CMN_LDO_M0_CFG_VREF_CTRL_FIELD 7:0
`define DDR_CMN_LDO_M0_CFG_VREF_CTRL_FIELD_WIDTH 8
`define DDR_CMN_LDO_M0_CFG_RANGE 13:0
`define DDR_CMN_LDO_M0_CFG_WIDTH 14
`define DDR_CMN_LDO_M0_CFG_ADR 32'h00000020
`define DDR_CMN_LDO_M0_CFG_POR 32'h00000000
`define DDR_CMN_LDO_M0_CFG_MSK 32'h00003FFF

// Word Address 0x00000024 : DDR_CMN_LDO_M1_CFG (RW)
`define DDR_CMN_LDO_M1_CFG_ATST_SEL_FIELD 12:10
`define DDR_CMN_LDO_M1_CFG_ATST_SEL_FIELD_WIDTH 3
`define DDR_CMN_LDO_M1_CFG_EN_FIELD 8
`define DDR_CMN_LDO_M1_CFG_EN_FIELD_WIDTH 1
`define DDR_CMN_LDO_M1_CFG_HIZ_FIELD 13
`define DDR_CMN_LDO_M1_CFG_HIZ_FIELD_WIDTH 1
`define DDR_CMN_LDO_M1_CFG_TRAN_ENH_EN_FIELD 9
`define DDR_CMN_LDO_M1_CFG_TRAN_ENH_EN_FIELD_WIDTH 1
`define DDR_CMN_LDO_M1_CFG_VREF_CTRL_FIELD 7:0
`define DDR_CMN_LDO_M1_CFG_VREF_CTRL_FIELD_WIDTH 8
`define DDR_CMN_LDO_M1_CFG_RANGE 13:0
`define DDR_CMN_LDO_M1_CFG_WIDTH 14
`define DDR_CMN_LDO_M1_CFG_ADR 32'h00000024
`define DDR_CMN_LDO_M1_CFG_POR 32'h00000000
`define DDR_CMN_LDO_M1_CFG_MSK 32'h00003FFF

// Word Address 0x00000028 : DDR_CMN_CLK_CTRL_CFG (RW)
`define DDR_CMN_CLK_CTRL_CFG_GFCM_EN_FIELD 3
`define DDR_CMN_CLK_CTRL_CFG_GFCM_EN_FIELD_WIDTH 1
`define DDR_CMN_CLK_CTRL_CFG_PLL0_DIV_CLK_BYP_FIELD 0
`define DDR_CMN_CLK_CTRL_CFG_PLL0_DIV_CLK_BYP_FIELD_WIDTH 1
`define DDR_CMN_CLK_CTRL_CFG_PLL0_DIV_CLK_EN_FIELD 2
`define DDR_CMN_CLK_CTRL_CFG_PLL0_DIV_CLK_EN_FIELD_WIDTH 1
`define DDR_CMN_CLK_CTRL_CFG_PLL0_DIV_CLK_RST_FIELD 1
`define DDR_CMN_CLK_CTRL_CFG_PLL0_DIV_CLK_RST_FIELD_WIDTH 1
`define DDR_CMN_CLK_CTRL_CFG_RANGE 3:0
`define DDR_CMN_CLK_CTRL_CFG_WIDTH 4
`define DDR_CMN_CLK_CTRL_CFG_ADR 32'h00000028
`define DDR_CMN_CLK_CTRL_CFG_POR 32'h00000002
`define DDR_CMN_CLK_CTRL_CFG_MSK 32'h0000000F

// Word Address 0x00000038 : DDR_CMN_PMON_ANA_CFG (RW)
`define DDR_CMN_PMON_ANA_CFG_NAND_EN_FIELD 0
`define DDR_CMN_PMON_ANA_CFG_NAND_EN_FIELD_WIDTH 1
`define DDR_CMN_PMON_ANA_CFG_NOR_EN_FIELD 1
`define DDR_CMN_PMON_ANA_CFG_NOR_EN_FIELD_WIDTH 1
`define DDR_CMN_PMON_ANA_CFG_RANGE 1:0
`define DDR_CMN_PMON_ANA_CFG_WIDTH 2
`define DDR_CMN_PMON_ANA_CFG_ADR 32'h00000038
`define DDR_CMN_PMON_ANA_CFG_POR 32'h00000000
`define DDR_CMN_PMON_ANA_CFG_MSK 32'h00000003

// Word Address 0x0000003C : DDR_CMN_PMON_DIG_CFG (RW)
`define DDR_CMN_PMON_DIG_CFG_INITWAIT_FIELD 7:0
`define DDR_CMN_PMON_DIG_CFG_INITWAIT_FIELD_WIDTH 8
`define DDR_CMN_PMON_DIG_CFG_REFCLK_RST_FIELD 8
`define DDR_CMN_PMON_DIG_CFG_REFCLK_RST_FIELD_WIDTH 1
`define DDR_CMN_PMON_DIG_CFG_RANGE 8:0
`define DDR_CMN_PMON_DIG_CFG_WIDTH 9
`define DDR_CMN_PMON_DIG_CFG_ADR 32'h0000003C
`define DDR_CMN_PMON_DIG_CFG_POR 32'h00000100
`define DDR_CMN_PMON_DIG_CFG_MSK 32'h000001FF

// Word Address 0x00000040 : DDR_CMN_PMON_DIG_NAND_CFG (RW)
`define DDR_CMN_PMON_DIG_NAND_CFG_COUNT_EN_FIELD 12
`define DDR_CMN_PMON_DIG_NAND_CFG_COUNT_EN_FIELD_WIDTH 1
`define DDR_CMN_PMON_DIG_NAND_CFG_REFCOUNT_FIELD 11:0
`define DDR_CMN_PMON_DIG_NAND_CFG_REFCOUNT_FIELD_WIDTH 12
`define DDR_CMN_PMON_DIG_NAND_CFG_RANGE 12:0
`define DDR_CMN_PMON_DIG_NAND_CFG_WIDTH 13
`define DDR_CMN_PMON_DIG_NAND_CFG_ADR 32'h00000040
`define DDR_CMN_PMON_DIG_NAND_CFG_POR 32'h00000000
`define DDR_CMN_PMON_DIG_NAND_CFG_MSK 32'h00001FFF

// Word Address 0x00000044 : DDR_CMN_PMON_DIG_NOR_CFG (RW)
`define DDR_CMN_PMON_DIG_NOR_CFG_COUNT_EN_FIELD 12
`define DDR_CMN_PMON_DIG_NOR_CFG_COUNT_EN_FIELD_WIDTH 1
`define DDR_CMN_PMON_DIG_NOR_CFG_REFCOUNT_FIELD 11:0
`define DDR_CMN_PMON_DIG_NOR_CFG_REFCOUNT_FIELD_WIDTH 12
`define DDR_CMN_PMON_DIG_NOR_CFG_RANGE 12:0
`define DDR_CMN_PMON_DIG_NOR_CFG_WIDTH 13
`define DDR_CMN_PMON_DIG_NOR_CFG_ADR 32'h00000044
`define DDR_CMN_PMON_DIG_NOR_CFG_POR 32'h00000000
`define DDR_CMN_PMON_DIG_NOR_CFG_MSK 32'h00001FFF

// Word Address 0x00000048 : DDR_CMN_PMON_NAND_STA (R)
`define DDR_CMN_PMON_NAND_STA_COUNT_FIELD 23:0
`define DDR_CMN_PMON_NAND_STA_COUNT_FIELD_WIDTH 24
`define DDR_CMN_PMON_NAND_STA_DONE_FIELD 24
`define DDR_CMN_PMON_NAND_STA_DONE_FIELD_WIDTH 1
`define DDR_CMN_PMON_NAND_STA_RANGE 24:0
`define DDR_CMN_PMON_NAND_STA_WIDTH 25
`define DDR_CMN_PMON_NAND_STA_ADR 32'h00000048
`define DDR_CMN_PMON_NAND_STA_POR 32'h00000000
`define DDR_CMN_PMON_NAND_STA_MSK 32'h01FFFFFF

// Word Address 0x0000004C : DDR_CMN_PMON_NOR_STA (R)
`define DDR_CMN_PMON_NOR_STA_COUNT_FIELD 23:0
`define DDR_CMN_PMON_NOR_STA_COUNT_FIELD_WIDTH 24
`define DDR_CMN_PMON_NOR_STA_DONE_FIELD 24
`define DDR_CMN_PMON_NOR_STA_DONE_FIELD_WIDTH 1
`define DDR_CMN_PMON_NOR_STA_RANGE 24:0
`define DDR_CMN_PMON_NOR_STA_WIDTH 25
`define DDR_CMN_PMON_NOR_STA_ADR 32'h0000004C
`define DDR_CMN_PMON_NOR_STA_POR 32'h00000000
`define DDR_CMN_PMON_NOR_STA_MSK 32'h01FFFFFF

// Word Address 0x00000050 : DDR_CMN_CLK_STA (R)
`define DDR_CMN_CLK_STA_GFCM0_CLKA_SEL_FIELD 0
`define DDR_CMN_CLK_STA_GFCM0_CLKA_SEL_FIELD_WIDTH 1
`define DDR_CMN_CLK_STA_GFCM0_CLKB_SEL_FIELD 1
`define DDR_CMN_CLK_STA_GFCM0_CLKB_SEL_FIELD_WIDTH 1
`define DDR_CMN_CLK_STA_GFCM1_CLKA_SEL_FIELD 2
`define DDR_CMN_CLK_STA_GFCM1_CLKA_SEL_FIELD_WIDTH 1
`define DDR_CMN_CLK_STA_GFCM1_CLKB_SEL_FIELD 3
`define DDR_CMN_CLK_STA_GFCM1_CLKB_SEL_FIELD_WIDTH 1
`define DDR_CMN_CLK_STA_RANGE 3:0
`define DDR_CMN_CLK_STA_WIDTH 4
`define DDR_CMN_CLK_STA_ADR 32'h00000050
`define DDR_CMN_CLK_STA_POR 32'h00000000
`define DDR_CMN_CLK_STA_MSK 32'h0000000F

// Word Address 0x00000054 : DDR_CMN_RSTN_CFG (RW)
`define DDR_CMN_RSTN_CFG_RSTN_BS_DIN_FIELD 3
`define DDR_CMN_RSTN_CFG_RSTN_BS_DIN_FIELD_WIDTH 1
`define DDR_CMN_RSTN_CFG_RSTN_BS_ENA_FIELD 4
`define DDR_CMN_RSTN_CFG_RSTN_BS_ENA_FIELD_WIDTH 1
`define DDR_CMN_RSTN_CFG_RSTN_LPBK_ENA_FIELD 2
`define DDR_CMN_RSTN_CFG_RSTN_LPBK_ENA_FIELD_WIDTH 1
`define DDR_CMN_RSTN_CFG_RSTN_OVR_SEL_FIELD 0
`define DDR_CMN_RSTN_CFG_RSTN_OVR_SEL_FIELD_WIDTH 1
`define DDR_CMN_RSTN_CFG_RSTN_OVR_VAL_FIELD 1
`define DDR_CMN_RSTN_CFG_RSTN_OVR_VAL_FIELD_WIDTH 1
`define DDR_CMN_RSTN_CFG_RANGE 4:0
`define DDR_CMN_RSTN_CFG_WIDTH 5
`define DDR_CMN_RSTN_CFG_ADR 32'h00000054
`define DDR_CMN_RSTN_CFG_POR 32'h00000000
`define DDR_CMN_RSTN_CFG_MSK 32'h0000001F

// Word Address 0x00000058 : DDR_CMN_RSTN_STA (R)
`define DDR_CMN_RSTN_STA_RSTN_LPBK_FIELD 0
`define DDR_CMN_RSTN_STA_RSTN_LPBK_FIELD_WIDTH 1
`define DDR_CMN_RSTN_STA_RANGE 0:0
`define DDR_CMN_RSTN_STA_WIDTH 1
`define DDR_CMN_RSTN_STA_ADR 32'h00000058
`define DDR_CMN_RSTN_STA_POR 32'h00000000
`define DDR_CMN_RSTN_STA_MSK 32'h00000001
