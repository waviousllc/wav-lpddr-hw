/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s001
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 15762
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_clkmux_diff_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_lib, Cell - wphy_clkmux_diff_wphy_clkmux_3to1_diff, View -
//schematic
// LAST TIME SAVED: Sep 17 21:04:57 2020
// NETLIST TIME: Oct 27 02:03:19 2020
`timescale 1ps / 1ps 




 

module wphy_clkmux_diff_wphy_clkmux_3to1_diff (out_c, out_t, vdda, vss, in01_c, in01_t, 
    in10_c, in10_t, in11_c, in11_t, s);

output  out_c, out_t;

inout  vdda, vss;

input  in01_c, in01_t, in10_c, in10_t, in11_c, in11_t;

input [1:0]  s;

// Buses in the design

wire  [1:0]  sb;

wire  [1:0]  s_buf;


wphy_clkmux_diff_INV_D2_GL16_LVT INV7 ( .in(s00b), .vss(vss), .out(s00), .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV5_1 ( .in(s[1]), .vss(vss), .out(sb[1]), 
    .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV5_0 ( .in(s[0]), .vss(vss), .out(sb[0]), 
    .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV6_1 ( .in(sb[1]), .vss(vss), .out(s_buf[1]), 
    .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV6_0 ( .in(sb[0]), .vss(vss), .out(s_buf[0]), 
    .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV4 ( .in(s01b), .vss(vss), .out(s01), .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV3 ( .in(s10b), .vss(vss), .out(s10), .vdd(vdda));

wphy_clkmux_diff_INV_D2_GL16_LVT INV2 ( .in(s11b), .vss(vss), .out(s11), .vdd(vdda));

wphy_clkmux_diff_INV_D16_GL16_LVT INV9 ( .in(yb_c), .vss(vss), .out(out_c), .vdd(vdda));

wphy_clkmux_diff_INV_D16_GL16_LVT INV8 ( .in(yb_t), .vss(vss), .out(out_t), .vdd(vdda));

wphy_clkmux_diff_NAND2_D1_GL16_LVT NAND3 ( .tielo(vss), .vdd(vdda), .y(s00b), .vss(vss), 
    .tiehi(vdda), .b(sb[0]), .a(sb[1]));

wphy_clkmux_diff_NAND2_D1_GL16_LVT NAND2 ( .tielo(vss), .vdd(vdda), .y(s10b), .vss(vss), 
    .tiehi(vdda), .b(sb[0]), .a(s_buf[1]));

wphy_clkmux_diff_NAND2_D1_GL16_LVT NAND1 ( .tielo(vss), .vdd(vdda), .y(s11b), .vss(vss), 
    .tiehi(vdda), .b(s_buf[0]), .a(s_buf[1]));

wphy_clkmux_diff_NAND2_D1_GL16_LVT NAND0 ( .tielo(vss), .vdd(vdda), .y(s01b), .vss(vss), 
    .tiehi(vdda), .b(s_buf[0]), .a(sb[1]));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT03_1 ( .out(mux_slw_cb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT03_0 ( .out(mux_slw_cb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT4_3 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT4_2 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT4_1 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT4_0 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT3_1 ( .out(mux_slw_tb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT3_0 ( .out(mux_slw_tb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT1_3 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT1_2 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT1_1 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT1_0 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT02_1 ( .out(mux_slw_cb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT02_0 ( .out(mux_slw_cb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_c), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT5_3 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT5_2 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT5_1 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT5_0 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT2_1 ( .out(mux_slw_tb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT2_0 ( .out(mux_slw_tb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT01_3 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT01_2 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT01_1 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_diff_INVT_D2_GL16_LVT INVT01_0 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_diff_PD_D1_GL16_LVT PD0 ( .vss(vss), .enb(s00), .y(yb_c));

wphy_clkmux_diff_PU_D1_GL16_LVT PU0 ( .vdd(vdda), .en(s00b), .y(yb_t));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_clkmux_diff, View -
//schematic
// LAST TIME SAVED: Sep 17 21:05:09 2020
// NETLIST TIME: Oct 27 02:03:19 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_clkmux_diff (d_ddrclk_c, d_ddrclk_t, d_qdrclk_c, 
    d_qdrclk_t,   d_ddrclk_sel, d_pi0, d_pi90, d_pi180, 
    d_pi270, d_qclk1_c, d_qclk1_t, d_qclk2_c, d_qclk2_t, d_qdrclk_sel, 
    d_rdqs_c, d_rdqs_t, d_wck_c, d_wck_t
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  d_ddrclk_c, d_ddrclk_t, d_qdrclk_c, d_qdrclk_t;



input  d_pi0, d_pi90, d_pi180, d_pi270, d_qclk1_c, d_qclk1_t, 
    d_qclk2_c, d_qclk2_t, d_rdqs_c, d_rdqs_t, d_wck_c, d_wck_t;

input [1:0]  d_ddrclk_sel;
input [1:0]  d_qdrclk_sel;

`ifdef SYNTHESIS
`else 

wphy_clkmux_diff_wphy_clkmux_3to1_diff MUX_QDR ( .vdda(vdda), .vss(vss), 
    .out_c(d_qdrclk_c), .out_t(d_qdrclk_t), .in01_c(d_qclk1_c), 
    .in01_t(d_qclk1_t), .in10_c(d_qclk2_c), .in10_t(d_qclk2_t), 
    .in11_c(d_pi270), .in11_t(d_pi90), .s(d_qdrclk_sel[1:0]));

wphy_clkmux_diff_wphy_clkmux_3to1_diff MUX_DDR ( .vdda(vdda), .vss(vss), 
    .out_c(d_ddrclk_c), .out_t(d_ddrclk_t), .in01_c(d_rdqs_c), 
    .in01_t(d_rdqs_t), .in10_c(d_wck_c), .in10_t(d_wck_t), 
    .in11_c(d_pi180), .in11_t(d_pi0), .s(d_ddrclk_sel[1:0]));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell - wphy_clkmux_diff_tb, View
//- schematic
// LAST TIME SAVED: Oct 26 23:43:56 2020
// NETLIST TIME: Oct 27 02:03:20 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_diff_PU_D1_GL16_LVT" "systemVerilog"


module wphy_clkmux_diff_PU_D1_GL16_LVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_diff_PD_D1_GL16_LVT" "systemVerilog"

module wphy_clkmux_diff_PD_D1_GL16_LVT( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_diff_INVT_D2_GL16_LVT" "systemVerilog"

module wphy_clkmux_diff_INVT_D2_GL16_LVT( in, out, en, enb 
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG



assign out = (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_diff_NAND2_D1_GL16_LVT" "systemVerilog"


module wphy_clkmux_diff_NAND2_D1_GL16_LVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_clkmux_diff_INV_D16_GL16_LVT" "systemVerilog"


module wphy_clkmux_diff_INV_D16_GL16_LVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_diff_INV_D2_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_clkmux_diff_INV_D2_GL16_LVT( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

    assign  out = ~in;

endmodule
`endif //SYNTHESIS
