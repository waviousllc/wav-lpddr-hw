/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 683
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_2to1_14g_rvt_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_lib, Cell - wphy_2to1_14g_rvt, View -
//schematic
// LAST TIME SAVED: Dec 30 13:10:56 2020
// NETLIST TIME: Jan 21 09:52:23 2021
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_2to1_14g_rvt (o_z,   i_clk, i_clk_b, i_dataf, 
    i_datar
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  o_z;



input  i_clk, i_clk_b, i_dataf, i_datar;

`ifdef SYNTHESIS
`else 

wphy_2to1_14g_rvt_wphy_2to1_lat_hz_rvt LA1 ( .vss(vss), .vdda(vdda), .d(i_datar), 
    .clkb(i_clk_b), .clk(i_clk), .q(o_z));

wphy_2to1_14g_rvt_wphy_2to1_lat_hz_rvt LA2 ( .vss(vss), .vdda(vdda), .d(net12), 
    .clkb(i_clk), .clk(i_clk_b), .q(o_z));

wphy_2to1_14g_rvt_LAT_D1_GL16_RVT LA0 ( .tielo(vss), .vss(vss), .vdd(vdda), .tiehi(vdda), 
    .d(i_dataf), .clkb(i_clk_b), .clk(i_clk), .q(net12));

`ifdef WPHY_ANA_TIMING

specify

  (i_clk   => o_z)   = 23;
  $setup(i_datar,posedge i_clk,30);
  //$hold(posedge i_clk,i_datar,-45);
  $setup(i_dataf,posedge i_clk,30);
  //$hold(posedge i_clk,i_dataf,-45);

endspecify

`endif

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell - wphy_2to1_14g_rvt_tb, View
//- schematic
// LAST TIME SAVED: Jan 21 09:29:22 2021
// NETLIST TIME: Jan 21 09:52:23 2021
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_2to1_14g_rvt_LAT_D1_GL16_RVT" "systemVerilog"

`timescale 1ps/1ps
module wphy_2to1_14g_rvt_LAT_D1_GL16_RVT( q, clk, clkb, d
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
);
 
  input clk;
  output q;  
  input d;
  input clkb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG


  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;

  assign q = (power_ok) ? 1'bz : 1'bx;
  
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ?
                           (clkb) ?
                                  (d===1'bx) ? $random : d
                                  : q
                           : 1'bx;

endmodule
//Verilog HDL for "wmx_d2d_serdes_lib", "wmx_LAT_D1_GL16_LVT_HZ" "functional"

`timescale 1ps/1ps
module wphy_2to1_14g_rvt_wphy_2to1_lat_hz_rvt ( q, vdda, vss, clk, clkb, d );

  output q;
  inout vdda;
  input d;
  input clk;
  input clkb;
  inout vss;

  reg q_int;
  reg q;
  wire polarity_ok = clk^clkb;
  wire pwr_ok = ~vss&vdda;
  initial begin
    q_int = $random;
  end

always @(*) begin
  if(clkb) begin
	q_int = (d === 1'bx) ? $random : d;
  end 
end 

always @(*) begin
#1	q = (polarity_ok&pwr_ok) ? (clk ? q_int : 1'bz) :1'bx;
end

endmodule
`endif //SYNTHESIS
