/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
****************************************************************************
*
* Module    : wav_mcutop_csr_defs.vh
* Date      : 2021-01-15
* Desciption: Autogenerated CSR block.
*
* $Id: wav_mcutop_csr_defs.vh,v 1.8 2021/01/15 19:26:39 schilukuri Exp $
*
****************************************************************************/

// Word Address 0x00000000 : WAV_MCUTOP_RSVD (RW)
`define WAV_MCUTOP_RSVD_RSVD_FIELD 31:0
`define WAV_MCUTOP_RSVD_RSVD_FIELD_WIDTH 32
`define WAV_MCUTOP_RSVD_RANGE 31:0
`define WAV_MCUTOP_RSVD_WIDTH 32
`define WAV_MCUTOP_RSVD_ADR 32'h00000000
`define WAV_MCUTOP_RSVD_POR 32'h00000000
`define WAV_MCUTOP_RSVD_MSK 32'hFFFFFFFF

// Word Address 0x00000004 : WAV_MCUTOP_CFG (RW)
`define WAV_MCUTOP_CFG_DEBUG_EN_FIELD 1
`define WAV_MCUTOP_CFG_DEBUG_EN_FIELD_WIDTH 1
`define WAV_MCUTOP_CFG_FETCH_EN_FIELD 0
`define WAV_MCUTOP_CFG_FETCH_EN_FIELD_WIDTH 1
`define WAV_MCUTOP_CFG_RANGE 1:0
`define WAV_MCUTOP_CFG_WIDTH 2
`define WAV_MCUTOP_CFG_ADR 32'h00000004
`define WAV_MCUTOP_CFG_POR 32'h00000000
`define WAV_MCUTOP_CFG_MSK 32'h00000003

// Word Address 0x00000008 : WAV_MCUTOP_STA (R)
`define WAV_MCUTOP_STA_RESERVED_FIELD 31:0
`define WAV_MCUTOP_STA_RESERVED_FIELD_WIDTH 32
`define WAV_MCUTOP_STA_RANGE 31:0
`define WAV_MCUTOP_STA_WIDTH 32
`define WAV_MCUTOP_STA_ADR 32'h00000008
`define WAV_MCUTOP_STA_POR 32'h00000000
`define WAV_MCUTOP_STA_MSK 32'hFFFFFFFF
