/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
****************************************************************************
*
* Module    : ddr_dfich_csr_defs.vh
* Date      : 2021-04-22
* Desciption: Autogenerated CSR block.
*
* $Id: ddr_dfich_csr_defs.vh,v 1.34 2021/04/23 22:16:10 mclovis Exp $
*
****************************************************************************/

// Word Address 0x00000000 : DDR_DFICH_TOP_1_CFG (RW)
`define DDR_DFICH_TOP_1_CFG_BUF_CLK_EN_FIELD 13
`define DDR_DFICH_TOP_1_CFG_BUF_CLK_EN_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_BUF_MODE_FIELD 12
`define DDR_DFICH_TOP_1_CFG_BUF_MODE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_CA_RDDATA_EN_FIELD 17
`define DDR_DFICH_TOP_1_CFG_CA_RDDATA_EN_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_DQBYTE_RDVALID_MASK_FIELD 31:28
`define DDR_DFICH_TOP_1_CFG_DQBYTE_RDVALID_MASK_FIELD_WIDTH 4
`define DDR_DFICH_TOP_1_CFG_RDATA_CLR_FIELD 8
`define DDR_DFICH_TOP_1_CFG_RDATA_CLR_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_RDATA_ENABLE_FIELD 9
`define DDR_DFICH_TOP_1_CFG_RDATA_ENABLE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_RDATA_UPDATE_FIELD 10
`define DDR_DFICH_TOP_1_CFG_RDATA_UPDATE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_RDOUT_EN_OVR_FIELD 19
`define DDR_DFICH_TOP_1_CFG_RDOUT_EN_OVR_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_RDOUT_EN_OVR_SEL_FIELD 18
`define DDR_DFICH_TOP_1_CFG_RDOUT_EN_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_TS_ENABLE_FIELD 0
`define DDR_DFICH_TOP_1_CFG_TS_ENABLE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_TS_RESET_FIELD 1
`define DDR_DFICH_TOP_1_CFG_TS_RESET_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_WCK_MODE_FIELD 16
`define DDR_DFICH_TOP_1_CFG_WCK_MODE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_WDATA_CLR_FIELD 4
`define DDR_DFICH_TOP_1_CFG_WDATA_CLR_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_WDATA_ENABLE_FIELD 6
`define DDR_DFICH_TOP_1_CFG_WDATA_ENABLE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_WDATA_HOLD_FIELD 5
`define DDR_DFICH_TOP_1_CFG_WDATA_HOLD_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_WDATA_UPDATE_FIELD 7
`define DDR_DFICH_TOP_1_CFG_WDATA_UPDATE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_1_CFG_RANGE 31:0
`define DDR_DFICH_TOP_1_CFG_WIDTH 32
`define DDR_DFICH_TOP_1_CFG_ADR 32'h00000000
`define DDR_DFICH_TOP_1_CFG_POR 32'h00002000
`define DDR_DFICH_TOP_1_CFG_MSK 32'hF00F37F3

// Word Address 0x00000004 : DDR_DFICH_TOP_2_CFG (RW)
`define DDR_DFICH_TOP_2_CFG_IG_LOAD_PTR_FIELD 1
`define DDR_DFICH_TOP_2_CFG_IG_LOAD_PTR_FIELD_WIDTH 1
`define DDR_DFICH_TOP_2_CFG_IG_LOOP_MODE_FIELD 0
`define DDR_DFICH_TOP_2_CFG_IG_LOOP_MODE_FIELD_WIDTH 1
`define DDR_DFICH_TOP_2_CFG_IG_NUM_LOOPS_FIELD 7:4
`define DDR_DFICH_TOP_2_CFG_IG_NUM_LOOPS_FIELD_WIDTH 4
`define DDR_DFICH_TOP_2_CFG_IG_START_PTR_FIELD 21:16
`define DDR_DFICH_TOP_2_CFG_IG_START_PTR_FIELD_WIDTH 6
`define DDR_DFICH_TOP_2_CFG_IG_STOP_PTR_FIELD 13:8
`define DDR_DFICH_TOP_2_CFG_IG_STOP_PTR_FIELD_WIDTH 6
`define DDR_DFICH_TOP_2_CFG_RANGE 21:0
`define DDR_DFICH_TOP_2_CFG_WIDTH 22
`define DDR_DFICH_TOP_2_CFG_ADR 32'h00000004
`define DDR_DFICH_TOP_2_CFG_POR 32'h00000010
`define DDR_DFICH_TOP_2_CFG_MSK 32'h003F3FF3

// Word Address 0x00000008 : DDR_DFICH_TOP_3_CFG (RW)
`define DDR_DFICH_TOP_3_CFG_TS_BRKPT_EN_FIELD 16
`define DDR_DFICH_TOP_3_CFG_TS_BRKPT_EN_FIELD_WIDTH 1
`define DDR_DFICH_TOP_3_CFG_TS_BRKPT_VAL_FIELD 15:0
`define DDR_DFICH_TOP_3_CFG_TS_BRKPT_VAL_FIELD_WIDTH 16
`define DDR_DFICH_TOP_3_CFG_RANGE 16:0
`define DDR_DFICH_TOP_3_CFG_WIDTH 17
`define DDR_DFICH_TOP_3_CFG_ADR 32'h00000008
`define DDR_DFICH_TOP_3_CFG_POR 32'h00000000
`define DDR_DFICH_TOP_3_CFG_MSK 32'h0001FFFF

// Word Address 0x0000000C : DDR_DFICH_TOP_STA (R)
`define DDR_DFICH_TOP_STA_EG_STATE_FIELD 5:4
`define DDR_DFICH_TOP_STA_EG_STATE_FIELD_WIDTH 2
`define DDR_DFICH_TOP_STA_EG_STATE_UPD_FIELD 6
`define DDR_DFICH_TOP_STA_EG_STATE_UPD_FIELD_WIDTH 1
`define DDR_DFICH_TOP_STA_IG_STATE_FIELD 1:0
`define DDR_DFICH_TOP_STA_IG_STATE_FIELD_WIDTH 2
`define DDR_DFICH_TOP_STA_IG_STATE_UPD_FIELD 2
`define DDR_DFICH_TOP_STA_IG_STATE_UPD_FIELD_WIDTH 1
`define DDR_DFICH_TOP_STA_RANGE 6:0
`define DDR_DFICH_TOP_STA_WIDTH 7
`define DDR_DFICH_TOP_STA_ADR 32'h0000000C
`define DDR_DFICH_TOP_STA_POR 32'h00000000
`define DDR_DFICH_TOP_STA_MSK 32'h00000077

// Word Address 0x00000010 : DDR_DFICH_IG_DATA_CFG (RW)
`define DDR_DFICH_IG_DATA_CFG_WDATA_FIELD 31:0
`define DDR_DFICH_IG_DATA_CFG_WDATA_FIELD_WIDTH 32
`define DDR_DFICH_IG_DATA_CFG_RANGE 31:0
`define DDR_DFICH_IG_DATA_CFG_WIDTH 32
`define DDR_DFICH_IG_DATA_CFG_ADR 32'h00000010
`define DDR_DFICH_IG_DATA_CFG_POR 32'h00000000
`define DDR_DFICH_IG_DATA_CFG_MSK 32'hFFFFFFFF

// Word Address 0x00000014 : DDR_DFICH_EG_DATA_STA (R)
`define DDR_DFICH_EG_DATA_STA_RDATA_FIELD 31:0
`define DDR_DFICH_EG_DATA_STA_RDATA_FIELD_WIDTH 32
`define DDR_DFICH_EG_DATA_STA_RANGE 31:0
`define DDR_DFICH_EG_DATA_STA_WIDTH 32
`define DDR_DFICH_EG_DATA_STA_ADR 32'h00000014
`define DDR_DFICH_EG_DATA_STA_POR 32'h00000000
`define DDR_DFICH_EG_DATA_STA_MSK 32'hFFFFFFFF

// Word Address 0x00000018 : DDR_DFICH_WRC_M0_CFG (RW)
`define DDR_DFICH_WRC_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WRC_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WRC_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WRC_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WRC_M0_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_WRC_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_WRC_M0_CFG_RANGE 15:0
`define DDR_DFICH_WRC_M0_CFG_WIDTH 16
`define DDR_DFICH_WRC_M0_CFG_ADR 32'h00000018
`define DDR_DFICH_WRC_M0_CFG_POR 32'h00005000
`define DDR_DFICH_WRC_M0_CFG_MSK 32'h0000F031

// Word Address 0x0000001C : DDR_DFICH_WRC_M1_CFG (RW)
`define DDR_DFICH_WRC_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WRC_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WRC_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WRC_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WRC_M1_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_WRC_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_WRC_M1_CFG_RANGE 15:0
`define DDR_DFICH_WRC_M1_CFG_WIDTH 16
`define DDR_DFICH_WRC_M1_CFG_ADR 32'h0000001C
`define DDR_DFICH_WRC_M1_CFG_POR 32'h00005000
`define DDR_DFICH_WRC_M1_CFG_MSK 32'h0000F031

// Word Address 0x00000020 : DDR_DFICH_WRCCTRL_M0_CFG (RW)
`define DDR_DFICH_WRCCTRL_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WRCCTRL_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WRCCTRL_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WRCCTRL_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WRCCTRL_M0_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_WRCCTRL_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_WRCCTRL_M0_CFG_RANGE 15:0
`define DDR_DFICH_WRCCTRL_M0_CFG_WIDTH 16
`define DDR_DFICH_WRCCTRL_M0_CFG_ADR 32'h00000020
`define DDR_DFICH_WRCCTRL_M0_CFG_POR 32'h00005000
`define DDR_DFICH_WRCCTRL_M0_CFG_MSK 32'h0000F031

// Word Address 0x00000024 : DDR_DFICH_WRCCTRL_M1_CFG (RW)
`define DDR_DFICH_WRCCTRL_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WRCCTRL_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WRCCTRL_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WRCCTRL_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WRCCTRL_M1_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_WRCCTRL_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_WRCCTRL_M1_CFG_RANGE 15:0
`define DDR_DFICH_WRCCTRL_M1_CFG_WIDTH 16
`define DDR_DFICH_WRCCTRL_M1_CFG_ADR 32'h00000024
`define DDR_DFICH_WRCCTRL_M1_CFG_POR 32'h00005000
`define DDR_DFICH_WRCCTRL_M1_CFG_MSK 32'h0000F031

// Word Address 0x00000028 : DDR_DFICH_CKCTRL_M0_CFG (RW)
`define DDR_DFICH_CKCTRL_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_CKCTRL_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_CKCTRL_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_CKCTRL_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_CKCTRL_M0_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_CKCTRL_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_CKCTRL_M0_CFG_RANGE 15:0
`define DDR_DFICH_CKCTRL_M0_CFG_WIDTH 16
`define DDR_DFICH_CKCTRL_M0_CFG_ADR 32'h00000028
`define DDR_DFICH_CKCTRL_M0_CFG_POR 32'h00005000
`define DDR_DFICH_CKCTRL_M0_CFG_MSK 32'h0000F031

// Word Address 0x0000002C : DDR_DFICH_CKCTRL_M1_CFG (RW)
`define DDR_DFICH_CKCTRL_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_CKCTRL_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_CKCTRL_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_CKCTRL_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_CKCTRL_M1_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_CKCTRL_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_CKCTRL_M1_CFG_RANGE 15:0
`define DDR_DFICH_CKCTRL_M1_CFG_WIDTH 16
`define DDR_DFICH_CKCTRL_M1_CFG_ADR 32'h0000002C
`define DDR_DFICH_CKCTRL_M1_CFG_POR 32'h00005000
`define DDR_DFICH_CKCTRL_M1_CFG_MSK 32'h0000F031

// Word Address 0x00000030 : DDR_DFICH_RDC_M0_CFG (RW)
`define DDR_DFICH_RDC_M0_CFG_GB_MODE_FIELD 3:0
`define DDR_DFICH_RDC_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_RDC_M0_CFG_RANGE 3:0
`define DDR_DFICH_RDC_M0_CFG_WIDTH 4
`define DDR_DFICH_RDC_M0_CFG_ADR 32'h00000030
`define DDR_DFICH_RDC_M0_CFG_POR 32'h00000006
`define DDR_DFICH_RDC_M0_CFG_MSK 32'h0000000F

// Word Address 0x00000034 : DDR_DFICH_RDC_M1_CFG (RW)
`define DDR_DFICH_RDC_M1_CFG_GB_MODE_FIELD 3:0
`define DDR_DFICH_RDC_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_RDC_M1_CFG_RANGE 3:0
`define DDR_DFICH_RDC_M1_CFG_WIDTH 4
`define DDR_DFICH_RDC_M1_CFG_ADR 32'h00000034
`define DDR_DFICH_RDC_M1_CFG_POR 32'h00000006
`define DDR_DFICH_RDC_M1_CFG_MSK 32'h0000000F

// Word Address 0x00000038 : DDR_DFICH_RCTRL_M0_CFG (RW)
`define DDR_DFICH_RCTRL_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_RCTRL_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_RCTRL_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_RCTRL_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_RCTRL_M0_CFG_POST_GB_FC_DLY_FIELD 6:4
`define DDR_DFICH_RCTRL_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 3
`define DDR_DFICH_RCTRL_M0_CFG_RANGE 15:0
`define DDR_DFICH_RCTRL_M0_CFG_WIDTH 16
`define DDR_DFICH_RCTRL_M0_CFG_ADR 32'h00000038
`define DDR_DFICH_RCTRL_M0_CFG_POR 32'h00005000
`define DDR_DFICH_RCTRL_M0_CFG_MSK 32'h0000F071

// Word Address 0x0000003C : DDR_DFICH_RCTRL_M1_CFG (RW)
`define DDR_DFICH_RCTRL_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_RCTRL_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_RCTRL_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_RCTRL_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_RCTRL_M1_CFG_POST_GB_FC_DLY_FIELD 6:4
`define DDR_DFICH_RCTRL_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 3
`define DDR_DFICH_RCTRL_M1_CFG_RANGE 15:0
`define DDR_DFICH_RCTRL_M1_CFG_WIDTH 16
`define DDR_DFICH_RCTRL_M1_CFG_ADR 32'h0000003C
`define DDR_DFICH_RCTRL_M1_CFG_POR 32'h00005000
`define DDR_DFICH_RCTRL_M1_CFG_MSK 32'h0000F071

// Word Address 0x00000040 : DDR_DFICH_WCTRL_M0_CFG (RW)
`define DDR_DFICH_WCTRL_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WCTRL_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WCTRL_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WCTRL_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WCTRL_M0_CFG_POST_GB_FC_DLY_FIELD 6:4
`define DDR_DFICH_WCTRL_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 3
`define DDR_DFICH_WCTRL_M0_CFG_RANGE 15:0
`define DDR_DFICH_WCTRL_M0_CFG_WIDTH 16
`define DDR_DFICH_WCTRL_M0_CFG_ADR 32'h00000040
`define DDR_DFICH_WCTRL_M0_CFG_POR 32'h00005000
`define DDR_DFICH_WCTRL_M0_CFG_MSK 32'h0000F071

// Word Address 0x00000044 : DDR_DFICH_WCTRL_M1_CFG (RW)
`define DDR_DFICH_WCTRL_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WCTRL_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WCTRL_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WCTRL_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WCTRL_M1_CFG_POST_GB_FC_DLY_FIELD 6:4
`define DDR_DFICH_WCTRL_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 3
`define DDR_DFICH_WCTRL_M1_CFG_RANGE 15:0
`define DDR_DFICH_WCTRL_M1_CFG_WIDTH 16
`define DDR_DFICH_WCTRL_M1_CFG_ADR 32'h00000044
`define DDR_DFICH_WCTRL_M1_CFG_POR 32'h00005000
`define DDR_DFICH_WCTRL_M1_CFG_MSK 32'h0000F071

// Word Address 0x00000048 : DDR_DFICH_WENCTRL_M0_CFG (RW)
`define DDR_DFICH_WENCTRL_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WENCTRL_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WENCTRL_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WENCTRL_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WENCTRL_M0_CFG_POST_GB_FC_DLY_FIELD 7:4
`define DDR_DFICH_WENCTRL_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 4
`define DDR_DFICH_WENCTRL_M0_CFG_RANGE 15:0
`define DDR_DFICH_WENCTRL_M0_CFG_WIDTH 16
`define DDR_DFICH_WENCTRL_M0_CFG_ADR 32'h00000048
`define DDR_DFICH_WENCTRL_M0_CFG_POR 32'h00005000
`define DDR_DFICH_WENCTRL_M0_CFG_MSK 32'h0000F0F1

// Word Address 0x0000004C : DDR_DFICH_WENCTRL_M1_CFG (RW)
`define DDR_DFICH_WENCTRL_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WENCTRL_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WENCTRL_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WENCTRL_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WENCTRL_M1_CFG_POST_GB_FC_DLY_FIELD 7:4
`define DDR_DFICH_WENCTRL_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 4
`define DDR_DFICH_WENCTRL_M1_CFG_RANGE 15:0
`define DDR_DFICH_WENCTRL_M1_CFG_WIDTH 16
`define DDR_DFICH_WENCTRL_M1_CFG_ADR 32'h0000004C
`define DDR_DFICH_WENCTRL_M1_CFG_POR 32'h00005000
`define DDR_DFICH_WENCTRL_M1_CFG_MSK 32'h0000F0F1

// Word Address 0x00000050 : DDR_DFICH_WCKCTRL_M0_CFG (RW)
`define DDR_DFICH_WCKCTRL_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WCKCTRL_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WCKCTRL_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WCKCTRL_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WCKCTRL_M0_CFG_POST_GB_FC_DLY_FIELD 6:4
`define DDR_DFICH_WCKCTRL_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 3
`define DDR_DFICH_WCKCTRL_M0_CFG_RANGE 15:0
`define DDR_DFICH_WCKCTRL_M0_CFG_WIDTH 16
`define DDR_DFICH_WCKCTRL_M0_CFG_ADR 32'h00000050
`define DDR_DFICH_WCKCTRL_M0_CFG_POR 32'h00005000
`define DDR_DFICH_WCKCTRL_M0_CFG_MSK 32'h0000F071

// Word Address 0x00000054 : DDR_DFICH_WCKCTRL_M1_CFG (RW)
`define DDR_DFICH_WCKCTRL_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WCKCTRL_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WCKCTRL_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WCKCTRL_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WCKCTRL_M1_CFG_POST_GB_FC_DLY_FIELD 6:4
`define DDR_DFICH_WCKCTRL_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 3
`define DDR_DFICH_WCKCTRL_M1_CFG_RANGE 15:0
`define DDR_DFICH_WCKCTRL_M1_CFG_WIDTH 16
`define DDR_DFICH_WCKCTRL_M1_CFG_ADR 32'h00000054
`define DDR_DFICH_WCKCTRL_M1_CFG_POR 32'h00005000
`define DDR_DFICH_WCKCTRL_M1_CFG_MSK 32'h0000F071

// Word Address 0x00000058 : DDR_DFICH_WRD_M0_CFG (RW)
`define DDR_DFICH_WRD_M0_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WRD_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WRD_M0_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WRD_M0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WRD_M0_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_WRD_M0_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_WRD_M0_CFG_RANGE 15:0
`define DDR_DFICH_WRD_M0_CFG_WIDTH 16
`define DDR_DFICH_WRD_M0_CFG_ADR 32'h00000058
`define DDR_DFICH_WRD_M0_CFG_POR 32'h00005000
`define DDR_DFICH_WRD_M0_CFG_MSK 32'h0000F031

// Word Address 0x0000005C : DDR_DFICH_WRD_M1_CFG (RW)
`define DDR_DFICH_WRD_M1_CFG_GB_MODE_FIELD 15:12
`define DDR_DFICH_WRD_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_WRD_M1_CFG_PIPE_EN_FIELD 0
`define DDR_DFICH_WRD_M1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_WRD_M1_CFG_POST_GB_FC_DLY_FIELD 5:4
`define DDR_DFICH_WRD_M1_CFG_POST_GB_FC_DLY_FIELD_WIDTH 2
`define DDR_DFICH_WRD_M1_CFG_RANGE 15:0
`define DDR_DFICH_WRD_M1_CFG_WIDTH 16
`define DDR_DFICH_WRD_M1_CFG_ADR 32'h0000005C
`define DDR_DFICH_WRD_M1_CFG_POR 32'h00005000
`define DDR_DFICH_WRD_M1_CFG_MSK 32'h0000F031

// Word Address 0x00000060 : DDR_DFICH_RDD_M0_CFG (RW)
`define DDR_DFICH_RDD_M0_CFG_GB_MODE_FIELD 3:0
`define DDR_DFICH_RDD_M0_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_RDD_M0_CFG_RANGE 3:0
`define DDR_DFICH_RDD_M0_CFG_WIDTH 4
`define DDR_DFICH_RDD_M0_CFG_ADR 32'h00000060
`define DDR_DFICH_RDD_M0_CFG_POR 32'h00000006
`define DDR_DFICH_RDD_M0_CFG_MSK 32'h0000000F

// Word Address 0x00000064 : DDR_DFICH_RDD_M1_CFG (RW)
`define DDR_DFICH_RDD_M1_CFG_GB_MODE_FIELD 3:0
`define DDR_DFICH_RDD_M1_CFG_GB_MODE_FIELD_WIDTH 4
`define DDR_DFICH_RDD_M1_CFG_RANGE 3:0
`define DDR_DFICH_RDD_M1_CFG_WIDTH 4
`define DDR_DFICH_RDD_M1_CFG_ADR 32'h00000064
`define DDR_DFICH_RDD_M1_CFG_POR 32'h00000006
`define DDR_DFICH_RDD_M1_CFG_MSK 32'h0000000F

// Word Address 0x00000068 : DDR_DFICH_CTRL0_M0_CFG (RW)
`define DDR_DFICH_CTRL0_M0_CFG_RD_INTF_PIPE_EN_FIELD 1
`define DDR_DFICH_CTRL0_M0_CFG_RD_INTF_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_CTRL0_M0_CFG_WR_INTF_PIPE_EN_FIELD 0
`define DDR_DFICH_CTRL0_M0_CFG_WR_INTF_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_CTRL0_M0_CFG_RANGE 1:0
`define DDR_DFICH_CTRL0_M0_CFG_WIDTH 2
`define DDR_DFICH_CTRL0_M0_CFG_ADR 32'h00000068
`define DDR_DFICH_CTRL0_M0_CFG_POR 32'h00000003
`define DDR_DFICH_CTRL0_M0_CFG_MSK 32'h00000003

// Word Address 0x0000006C : DDR_DFICH_CTRL0_M1_CFG (RW)
`define DDR_DFICH_CTRL0_M1_CFG_RD_INTF_PIPE_EN_FIELD 1
`define DDR_DFICH_CTRL0_M1_CFG_RD_INTF_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_CTRL0_M1_CFG_WR_INTF_PIPE_EN_FIELD 0
`define DDR_DFICH_CTRL0_M1_CFG_WR_INTF_PIPE_EN_FIELD_WIDTH 1
`define DDR_DFICH_CTRL0_M1_CFG_RANGE 1:0
`define DDR_DFICH_CTRL0_M1_CFG_WIDTH 2
`define DDR_DFICH_CTRL0_M1_CFG_ADR 32'h0000006C
`define DDR_DFICH_CTRL0_M1_CFG_POR 32'h00000003
`define DDR_DFICH_CTRL0_M1_CFG_MSK 32'h00000003

// Word Address 0x00000070 : DDR_DFICH_CTRL1_M0_CFG (RW)
`define DDR_DFICH_CTRL1_M0_CFG_CA_TRAFFIC_OVR_FIELD 6
`define DDR_DFICH_CTRL1_M0_CFG_CA_TRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_CA_TRAFFIC_OVR_SEL_FIELD 2
`define DDR_DFICH_CTRL1_M0_CFG_CA_TRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_CK_TRAFFIC_OVR_FIELD 7
`define DDR_DFICH_CTRL1_M0_CFG_CK_TRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_CK_TRAFFIC_OVR_SEL_FIELD 3
`define DDR_DFICH_CTRL1_M0_CFG_CK_TRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_DQS_WRTRAFFIC_OVR_FIELD 5
`define DDR_DFICH_CTRL1_M0_CFG_DQS_WRTRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_DQS_WRTRAFFIC_OVR_SEL_FIELD 1
`define DDR_DFICH_CTRL1_M0_CFG_DQS_WRTRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_DQ_RDTRAFFIC_OVR_FIELD 9
`define DDR_DFICH_CTRL1_M0_CFG_DQ_RDTRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_DQ_RDTRAFFIC_OVR_SEL_FIELD 8
`define DDR_DFICH_CTRL1_M0_CFG_DQ_RDTRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_DQ_WRTRAFFIC_OVR_FIELD 4
`define DDR_DFICH_CTRL1_M0_CFG_DQ_WRTRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_DQ_WRTRAFFIC_OVR_SEL_FIELD 0
`define DDR_DFICH_CTRL1_M0_CFG_DQ_WRTRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M0_CFG_RANGE 9:0
`define DDR_DFICH_CTRL1_M0_CFG_WIDTH 10
`define DDR_DFICH_CTRL1_M0_CFG_ADR 32'h00000070
`define DDR_DFICH_CTRL1_M0_CFG_POR 32'h000000FF
`define DDR_DFICH_CTRL1_M0_CFG_MSK 32'h000003FF

// Word Address 0x00000074 : DDR_DFICH_CTRL1_M1_CFG (RW)
`define DDR_DFICH_CTRL1_M1_CFG_CA_TRAFFIC_OVR_FIELD 6
`define DDR_DFICH_CTRL1_M1_CFG_CA_TRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_CA_TRAFFIC_OVR_SEL_FIELD 2
`define DDR_DFICH_CTRL1_M1_CFG_CA_TRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_CK_TRAFFIC_OVR_FIELD 7
`define DDR_DFICH_CTRL1_M1_CFG_CK_TRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_CK_TRAFFIC_OVR_SEL_FIELD 3
`define DDR_DFICH_CTRL1_M1_CFG_CK_TRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_DQS_WRTRAFFIC_OVR_FIELD 5
`define DDR_DFICH_CTRL1_M1_CFG_DQS_WRTRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_DQS_WRTRAFFIC_OVR_SEL_FIELD 1
`define DDR_DFICH_CTRL1_M1_CFG_DQS_WRTRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_DQ_RDTRAFFIC_OVR_FIELD 9
`define DDR_DFICH_CTRL1_M1_CFG_DQ_RDTRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_DQ_RDTRAFFIC_OVR_SEL_FIELD 8
`define DDR_DFICH_CTRL1_M1_CFG_DQ_RDTRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_DQ_WRTRAFFIC_OVR_FIELD 4
`define DDR_DFICH_CTRL1_M1_CFG_DQ_WRTRAFFIC_OVR_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_DQ_WRTRAFFIC_OVR_SEL_FIELD 0
`define DDR_DFICH_CTRL1_M1_CFG_DQ_WRTRAFFIC_OVR_SEL_FIELD_WIDTH 1
`define DDR_DFICH_CTRL1_M1_CFG_RANGE 9:0
`define DDR_DFICH_CTRL1_M1_CFG_WIDTH 10
`define DDR_DFICH_CTRL1_M1_CFG_ADR 32'h00000074
`define DDR_DFICH_CTRL1_M1_CFG_POR 32'h000000FF
`define DDR_DFICH_CTRL1_M1_CFG_MSK 32'h000003FF

// Word Address 0x00000078 : DDR_DFICH_CTRL2_M0_CFG (RW)
`define DDR_DFICH_CTRL2_M0_CFG_CA_CLK_EN_PULSE_EXT_FIELD 11:8
`define DDR_DFICH_CTRL2_M0_CFG_CA_CLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M0_CFG_CK_CLK_EN_PULSE_EXT_FIELD 15:12
`define DDR_DFICH_CTRL2_M0_CFG_CK_CLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M0_CFG_DQS_WRCLK_EN_PULSE_EXT_FIELD 7:4
`define DDR_DFICH_CTRL2_M0_CFG_DQS_WRCLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M0_CFG_DQ_WRCLK_EN_PULSE_EXT_FIELD 3:0
`define DDR_DFICH_CTRL2_M0_CFG_DQ_WRCLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M0_CFG_RDCLK_EN_PULSE_EXT_FIELD 19:16
`define DDR_DFICH_CTRL2_M0_CFG_RDCLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M0_CFG_RANGE 19:0
`define DDR_DFICH_CTRL2_M0_CFG_WIDTH 20
`define DDR_DFICH_CTRL2_M0_CFG_ADR 32'h00000078
`define DDR_DFICH_CTRL2_M0_CFG_POR 32'h000F0033
`define DDR_DFICH_CTRL2_M0_CFG_MSK 32'h000FFFFF

// Word Address 0x0000007C : DDR_DFICH_CTRL2_M1_CFG (RW)
`define DDR_DFICH_CTRL2_M1_CFG_CA_CLK_EN_PULSE_EXT_FIELD 11:8
`define DDR_DFICH_CTRL2_M1_CFG_CA_CLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M1_CFG_CK_CLK_EN_PULSE_EXT_FIELD 15:12
`define DDR_DFICH_CTRL2_M1_CFG_CK_CLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M1_CFG_DQS_WRCLK_EN_PULSE_EXT_FIELD 7:4
`define DDR_DFICH_CTRL2_M1_CFG_DQS_WRCLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M1_CFG_DQ_WRCLK_EN_PULSE_EXT_FIELD 3:0
`define DDR_DFICH_CTRL2_M1_CFG_DQ_WRCLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M1_CFG_RDCLK_EN_PULSE_EXT_FIELD 19:16
`define DDR_DFICH_CTRL2_M1_CFG_RDCLK_EN_PULSE_EXT_FIELD_WIDTH 4
`define DDR_DFICH_CTRL2_M1_CFG_RANGE 19:0
`define DDR_DFICH_CTRL2_M1_CFG_WIDTH 20
`define DDR_DFICH_CTRL2_M1_CFG_ADR 32'h0000007C
`define DDR_DFICH_CTRL2_M1_CFG_POR 32'h000F0033
`define DDR_DFICH_CTRL2_M1_CFG_MSK 32'h000FFFFF

// Word Address 0x00000080 : DDR_DFICH_CTRL3_M0_CFG (RW)
`define DDR_DFICH_CTRL3_M0_CFG_WRD_CS_PHASE_EXT_FIELD 5:0
`define DDR_DFICH_CTRL3_M0_CFG_WRD_CS_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL3_M0_CFG_WRD_EN_PHASE_EXT_FIELD 13:8
`define DDR_DFICH_CTRL3_M0_CFG_WRD_EN_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL3_M0_CFG_WRD_OE_PHASE_EXT_FIELD 21:16
`define DDR_DFICH_CTRL3_M0_CFG_WRD_OE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL3_M0_CFG_RANGE 21:0
`define DDR_DFICH_CTRL3_M0_CFG_WIDTH 22
`define DDR_DFICH_CTRL3_M0_CFG_ADR 32'h00000080
`define DDR_DFICH_CTRL3_M0_CFG_POR 32'h00020200
`define DDR_DFICH_CTRL3_M0_CFG_MSK 32'h003F3F3F

// Word Address 0x00000084 : DDR_DFICH_CTRL3_M1_CFG (RW)
`define DDR_DFICH_CTRL3_M1_CFG_WRD_CS_PHASE_EXT_FIELD 5:0
`define DDR_DFICH_CTRL3_M1_CFG_WRD_CS_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL3_M1_CFG_WRD_EN_PHASE_EXT_FIELD 13:8
`define DDR_DFICH_CTRL3_M1_CFG_WRD_EN_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL3_M1_CFG_WRD_OE_PHASE_EXT_FIELD 21:16
`define DDR_DFICH_CTRL3_M1_CFG_WRD_OE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL3_M1_CFG_RANGE 21:0
`define DDR_DFICH_CTRL3_M1_CFG_WIDTH 22
`define DDR_DFICH_CTRL3_M1_CFG_ADR 32'h00000084
`define DDR_DFICH_CTRL3_M1_CFG_POR 32'h00020200
`define DDR_DFICH_CTRL3_M1_CFG_MSK 32'h003F3F3F

// Word Address 0x00000088 : DDR_DFICH_CTRL4_M0_CFG (RW)
`define DDR_DFICH_CTRL4_M0_CFG_WCK_CS_PHASE_EXT_FIELD 13:8
`define DDR_DFICH_CTRL4_M0_CFG_WCK_CS_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL4_M0_CFG_WCK_OE_PHASE_EXT_FIELD 5:0
`define DDR_DFICH_CTRL4_M0_CFG_WCK_OE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL4_M0_CFG_RANGE 13:0
`define DDR_DFICH_CTRL4_M0_CFG_WIDTH 14
`define DDR_DFICH_CTRL4_M0_CFG_ADR 32'h00000088
`define DDR_DFICH_CTRL4_M0_CFG_POR 32'h00000002
`define DDR_DFICH_CTRL4_M0_CFG_MSK 32'h00003F3F

// Word Address 0x0000008C : DDR_DFICH_CTRL4_M1_CFG (RW)
`define DDR_DFICH_CTRL4_M1_CFG_WCK_CS_PHASE_EXT_FIELD 13:8
`define DDR_DFICH_CTRL4_M1_CFG_WCK_CS_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL4_M1_CFG_WCK_OE_PHASE_EXT_FIELD 5:0
`define DDR_DFICH_CTRL4_M1_CFG_WCK_OE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL4_M1_CFG_RANGE 13:0
`define DDR_DFICH_CTRL4_M1_CFG_WIDTH 14
`define DDR_DFICH_CTRL4_M1_CFG_ADR 32'h0000008C
`define DDR_DFICH_CTRL4_M1_CFG_POR 32'h00000002
`define DDR_DFICH_CTRL4_M1_CFG_MSK 32'h00003F3F

// Word Address 0x00000090 : DDR_DFICH_CTRL5_M0_CFG (RW)
`define DDR_DFICH_CTRL5_M0_CFG_IE_PHASE_EXT_FIELD 13:8
`define DDR_DFICH_CTRL5_M0_CFG_IE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M0_CFG_RCS_PHASE_EXT_FIELD 5:0
`define DDR_DFICH_CTRL5_M0_CFG_RCS_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M0_CFG_REN_PHASE_EXT_FIELD 29:24
`define DDR_DFICH_CTRL5_M0_CFG_REN_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M0_CFG_RE_PHASE_EXT_FIELD 21:16
`define DDR_DFICH_CTRL5_M0_CFG_RE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M0_CFG_RANGE 29:0
`define DDR_DFICH_CTRL5_M0_CFG_WIDTH 30
`define DDR_DFICH_CTRL5_M0_CFG_ADR 32'h00000090
`define DDR_DFICH_CTRL5_M0_CFG_POR 32'h00000000
`define DDR_DFICH_CTRL5_M0_CFG_MSK 32'h3F3F3F3F

// Word Address 0x00000094 : DDR_DFICH_CTRL5_M1_CFG (RW)
`define DDR_DFICH_CTRL5_M1_CFG_IE_PHASE_EXT_FIELD 13:8
`define DDR_DFICH_CTRL5_M1_CFG_IE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M1_CFG_RCS_PHASE_EXT_FIELD 5:0
`define DDR_DFICH_CTRL5_M1_CFG_RCS_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M1_CFG_REN_PHASE_EXT_FIELD 29:24
`define DDR_DFICH_CTRL5_M1_CFG_REN_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M1_CFG_RE_PHASE_EXT_FIELD 21:16
`define DDR_DFICH_CTRL5_M1_CFG_RE_PHASE_EXT_FIELD_WIDTH 6
`define DDR_DFICH_CTRL5_M1_CFG_RANGE 29:0
`define DDR_DFICH_CTRL5_M1_CFG_WIDTH 30
`define DDR_DFICH_CTRL5_M1_CFG_ADR 32'h00000094
`define DDR_DFICH_CTRL5_M1_CFG_POR 32'h00000000
`define DDR_DFICH_CTRL5_M1_CFG_MSK 32'h3F3F3F3F
