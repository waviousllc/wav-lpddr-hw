/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 37506
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_gfcm_lvt_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_lib, Cell - wphy_gfcm_lvt, View -
//schematic
// LAST TIME SAVED: Oct 26 15:31:23 2020
// NETLIST TIME: Nov  3 00:04:19 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_gfcm_lvt (o_clk0, o_clk180,   clk_sel, ena, 
    i_clka0, i_clka180, i_clkb0, i_clkb180
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  o_clk0, o_clk180;



input  clk_sel, ena, i_clka0, i_clka180, i_clkb0, i_clkb180;

`ifdef SYNTHESIS
`else 

wphy_gfcm_lvt_INV_D2_GL16_LVT INV2 ( .in(enb), .vss(vss), .out(en), .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV19 ( .in(pu_en), .vss(vss), .out(pd_enb), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV1 ( .in(clk_sel), .vss(vss), .out(clk_selb), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV16 ( .in(en_b), .vss(vss), .out(enb_b), .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV15_1 ( .in(net050), .vss(vss), .out(clkb180), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV15_0 ( .in(net050), .vss(vss), .out(clkb180), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV14_1 ( .in(net034), .vss(vss), .out(clkb0), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV14_0 ( .in(net034), .vss(vss), .out(clkb0), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV13 ( .in(i_clkb0), .vss(vss), .out(net034), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV12 ( .in(i_clkb180), .vss(vss), .out(net050), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV11_1 ( .in(net049), .vss(vss), .out(clka180), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV11_0 ( .in(net049), .vss(vss), .out(clka180), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV8 ( .in(i_clka0), .vss(vss), .out(net019), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT I1 ( .in(net5), .vss(vss), .out(net038), .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV0 ( .in(net2), .vss(vss), .out(net09), .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV3 ( .in(en_a), .vss(vss), .out(enb_a), .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV7 ( .in(net035), .vss(vss), .out(o_clk180), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV6 ( .in(net036), .vss(vss), .out(o_clk0), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV20 ( .in(ena), .vss(vss), .out(enb), .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV9_1 ( .in(net019), .vss(vss), .out(clka0), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV9_0 ( .in(net019), .vss(vss), .out(clka0), 
    .vdd(vdda));

wphy_gfcm_lvt_INV_D2_GL16_LVT INV10 ( .in(i_clka180), .vss(vss), .out(net049), 
    .vdd(vdda));

wphy_gfcm_lvt_INVT_D2_GL16_LVT INVT0 ( .out(net036), .en(en_a), .enb(enb_a), 
    .vss(vss), .in(clka0), .vdd(vdda));

wphy_gfcm_lvt_INVT_D2_GL16_LVT INVT5 ( .out(net035), .en(en_a), .enb(enb_a), 
    .vss(vss), .in(clka180), .vdd(vdda));

wphy_gfcm_lvt_INVT_D2_GL16_LVT INVT4 ( .out(net035), .en(en_b), .enb(enb_b), 
    .vss(vss), .in(clkb180), .vdd(vdda));

wphy_gfcm_lvt_INVT_D2_GL16_LVT INVT3 ( .out(net036), .en(en_b), .enb(enb_b), 
    .vss(vss), .in(clkb0), .vdd(vdda));

wphy_gfcm_lvt_NOR2_D1_GL16_LVT NOR0 ( .tielo(vss), .tiehi(vdda), .y(sel_clkb), 
    .vss(vss), .vdd(vdda), .b(enb), .a(clk_selb));

wphy_gfcm_lvt_NOR2_D1_GL16_LVT NOR1 ( .tielo(vss), .tiehi(vdda), .y(sel_cala), 
    .vss(vss), .vdd(vdda), .b(enb), .a(sel_clkb));

wphy_gfcm_lvt_LATRES_D1_GL16_LVT LA0 ( .tielo(vss), .tiehi(vdda), .vss(vss), 
    .vdd(vdda), .rstb(en), .d(net09), .clkb(clkb180), .clk(clkb0), 
    .q(en_b));

wphy_gfcm_lvt_LATRES_D1_GL16_LVT LA00 ( .tielo(vss), .tiehi(vdda), .vss(vss), 
    .vdd(vdda), .rstb(en), .d(net038), .clkb(clka180), .clk(clka0), 
    .q(en_a));

wphy_gfcm_lvt_PU_D1_GL16_LVT PU0 ( .vdd(vdda), .en(pu_en), .y(net036));

wphy_gfcm_lvt_PD_D1_GL16_LVT PD0 ( .vss(vss), .enb(pd_enb), .y(net035));

wphy_gfcm_lvt_NAND2_D1_GL16_LVT NAND2 ( .tielo(vss), .vdd(vdda), .y(pu_en), 
    .vss(vss), .tiehi(vdda), .b(enb_b), .a(enb_a));

wphy_gfcm_lvt_NAND2_D1_GL16_LVT NAND1 ( .tielo(vss), .vdd(vdda), .y(net1), .vss(vss), 
    .tiehi(vdda), .b(net5), .a(sel_clkb));

wphy_gfcm_lvt_NAND2_D1_GL16_LVT NAND0 ( .tielo(vss), .vdd(vdda), .y(net4), .vss(vss), 
    .tiehi(vdda), .b(net2), .a(sel_cala));

wphy_gfcm_lvt_LATSET_D1_GL16_LVT LA1 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net6), .clkb(clka180), .clk(clka0), .q(net023));

wphy_gfcm_lvt_LATSET_D1_GL16_LVT LA4 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net3), .clkb(clkb180), .clk(clkb0), .q(net022));

wphy_gfcm_lvt_LATSET_D1_GL16_LVT LA2 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net023), .clkb(clka0), .clk(clka180), .q(net5));

wphy_gfcm_lvt_LATSET_D1_GL16_LVT LA3 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net022), .clkb(clkb0), .clk(clkb180), .q(net2));

wphy_gfcm_lvt_FFSET_D1_GL16_LVT FF0 ( .prst(enb), .prstb(en), .tielo(vss), .vss(vss), 
    .vdd(vdda), .tiehi(vdda), .d(net1), .clkb(clkb180), .clk(clkb0), 
    .q(net3));

wphy_gfcm_lvt_FFSET_D1_GL16_LVT FF1 ( .prst(enb), .prstb(en), .tielo(vss), .vss(vss), 
    .vdd(vdda), .tiehi(vdda), .d(net4), .clkb(clka180), .clk(clka0), 
    .q(net6));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell - wphy_gfcm_lvt_tb, View -
//schematic
// LAST TIME SAVED: Nov  2 23:58:10 2020
// NETLIST TIME: Nov  3 00:04:19 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_FFSET_D1_GL16_LVT" "systemVerilog"


module wphy_gfcm_lvt_FFSET_D1_GL16_LVT ( q, clk, clkb, d, prst, prstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input clk;
  input prst;
  input prstb;
  output q;
  input d;
  input clkb;   
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;

  initial  begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  initial  begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  reg q;

  initial begin
    q = $random;
  end

  always @(posedge clk or posedge prst) begin
   if(prst) begin
       q <= 1'b1;
    end else begin
       q <= d;
    end
  end

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_gfcm_lvt_LATSET_D1_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_gfcm_lvt_LATSET_D1_GL16_LVT ( q, clk, clkb, d, set
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo 
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  output q;
  input set;
  input d;
  input clk;
  input clkb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

assign #1  q = polarity_ok ? 
                           (set) ? 
                                 1'b1 
                                 : (clkb) ? 
                                          (d===1'bx) ? $random : d
                                          : q 
                           : 1'bx;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_NAND2_D1_GL16_LVT" "systemVerilog"


module wphy_gfcm_lvt_NAND2_D1_GL16_LVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_PD_D1_GL16_LVT" "systemVerilog"

module wphy_gfcm_lvt_PD_D1_GL16_LVT( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_PU_D1_GL16_LVT" "systemVerilog"


module wphy_gfcm_lvt_PU_D1_GL16_LVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_gfcm_lvt_LATRES_D1_GL16_LVT" "systemVerilog"


`timescale 1ps/1ps
module wphy_gfcm_lvt_LATRES_D1_GL16_LVT( q, clk, clkb, d, rstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo 
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PGL
);

  input clk;
  output q;
  input d;
  input clkb;
  input rstb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ? 
                           (~rstb) ? 
                                 1'b0 
                                 : (clkb) ? 
                                          (d===1'bx) ? $random : d&rstb
                                          : q 
                           : 1'bx;

endmodule

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_NOR2_D1_GL16_LVT" "systemVerilog"


module wphy_gfcm_lvt_NOR2_D1_GL16_LVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_INVT_D2_GL16_LVT" "systemVerilog"

module wphy_gfcm_lvt_INVT_D2_GL16_LVT( in, out, en, enb 
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG



assign out = (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_gfcm_lvt_INV_D2_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_gfcm_lvt_INV_D2_GL16_LVT( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

    assign  out = ~in;

endmodule
`endif //SYNTHESIS
