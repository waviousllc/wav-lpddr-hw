/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 35526
// Design library name: wphy_gf12lp_lp4x5_sim_lib
// Design cell name: wphy_lp4x5_cmn_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_wphy_lp4x5_cke_drvr_w_lpbk,
//View - schematic
// LAST TIME SAVED: Dec 14 16:29:59 2020
// NETLIST TIME: Jan 17 22:00:25 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_wphy_lp4x5_cke_drvr_w_lpbk (d_lpbk_out, pad_cke_out, vdda, 
    vdda1p2, vss, d_bs_din, d_bs_ena, d_in_c, d_lpbk_ena, d_ovrd, 
    d_ovrd_val, freeze_n_hv);

output  d_lpbk_out;

inout  pad_cke_out, vdda, vdda1p2, vss;

input  d_bs_din, d_bs_ena, d_in_c, d_lpbk_ena, d_ovrd_val, freeze_n_hv;

input [2:0]  d_ovrd;


wphy_lp4x5_cmn_MUXT2_D2_GL16_RVT MUX1 ( .vss(vss), .sb(bs_enb), .s(bs_ena), 
    .b(d_bs_din), .a(d_ovrd_val), .yb(ovrd_b_input), .vdd(vdda));

wphy_lp4x5_cmn_MUXT2_D2_GL16_RVT MUX0 ( .vss(vss), .sb(ovrdORbs), .s(ovrdNORbs), 
    .b(d_in_c), .a(ovrd_b_input), .yb(in_t), .vdd(vdda));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV3 ( .in(ovrdNORbs), .vss(vss), .out(ovrdORbs), 
    .vdd(vdda));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV6 ( .in(d_bs_ena), .vss(vss), .out(bs_enb), 
    .vdd(vdda));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV7 ( .in(bs_enb), .vss(vss), .out(bs_ena), 
    .vdd(vdda));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0 ( .in(ovrd_b), .vss(vss), .out(ovrd), .vdd(vdda));

wphy_lp4x5_cmn_NOR2_D1_GL16_LVT NOR1 ( .tielo(vss), .tiehi(vdda), .y(ovrdNORbs), 
    .vss(vss), .vdd(vdda), .b(bs_ena), .a(ovrd));

wphy_lp4x5_cmn_wphy_lp4x5_cke_drv_core DRV ( .vdda1p2(vdda1p2), .out_h(pad_cke_out), 
    .inb_h(inb_h), .vss(vss));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2 ( .vdda1p2(vdda), .in(net014), .vss(vss), 
    .out(d_lpbk_out));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0 ( .freezeb_hv(freeze_n_hv), 
    .outn(lpbk_enb_h), .in(d_lpbk_ena), .outp(lpbk_ena_h), 
    .vdda1p8(vdda1p2), .vdd(vdda), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LS0 ( .freezeb_hv(freeze_n_hv), .outn(inb_h), 
    .in(in_t), .outp(net015), .vdda1p8(vdda1p2), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_NOR3_D1_GL16_RVT NOR0 ( .vdd(vdda), .c(d_ovrd[0]), .y(ovrd_b), 
    .vss(vss), .b(d_ovrd[1]), .a(d_ovrd[2]));

wphy_lp4x5_cmn_cdm SEC_ESD1 ( .pad(pad_cke_out), .vdd(vdda1p2), .vss(vss), 
    .out(rxin_h));

wphy_lp4x5_cmn_hbm PRIM_ESD0_1 ( .vss(vss), .vdd(vdda1p2), .pad(pad_cke_out));

wphy_lp4x5_cmn_hbm PRIM_ESD0_0 ( .vss(vss), .vdd(vdda1p2), .pad(pad_cke_out));

wphy_lp4x5_cmn_NAND2_D1_GL150_EGU NAND0 ( .y(net014), .vss(vss), .vdda1p2(vdda1p2), 
    .b(lpbk_ena_h), .a(rxin_h));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_wphy_lp4x5_drv_240, View -
//schematic
// LAST TIME SAVED: Nov 30 15:42:35 2020
// NETLIST TIME: Jan 17 22:00:26 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_wphy_lp4x5_drv_240 (drv_out, vddq, vss, en_dn, en_up, inb_n, 
    inb_p, ncal, pcal);

output  drv_out;

inout  vddq, vss;

input  en_dn, en_up, inb_n, inb_p;

input [5:0]  pcal;
input [4:0]  ncal;

// Buses in the design

wire  [5:0]  nbb;

wire  [6:0]  p1;

wire  [6:0]  pb;

wire  [4:0]  net022;

wire  [6:0]  p;

wire  [5:0]  calp;

wire  [4:0]  dn_code;

wire  [5:0]  net023;

wire  [4:0]  caln;

wire  [5:0]  n1;

wire  [5:0]  n;

wire  [5:0]  up_code;


wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_240n I4 ( .out(drv_out), .dn_code(dn_code), 
    .dn_fix(n_fix), .vss(vss));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_6 ( .tiehi(vddq), .tielo(vss), .in(pb[6]), 
    .vss(vss), .out(p1[6]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_5 ( .tiehi(vddq), .tielo(vss), .in(pb[5]), 
    .vss(vss), .out(p1[5]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_4 ( .tiehi(vddq), .tielo(vss), .in(pb[4]), 
    .vss(vss), .out(p1[4]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_3 ( .tiehi(vddq), .tielo(vss), .in(pb[3]), 
    .vss(vss), .out(p1[3]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_2 ( .tiehi(vddq), .tielo(vss), .in(pb[2]), 
    .vss(vss), .out(p1[2]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_1 ( .tiehi(vddq), .tielo(vss), .in(pb[1]), 
    .vss(vss), .out(p1[1]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D1_GL16_SLVT INV1_0 ( .tiehi(vddq), .tielo(vss), .in(pb[0]), 
    .vss(vss), .out(p1[0]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV5_1 ( .in(p1[6]), .vss(vss), .out(p[6]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV5_0 ( .in(p1[5]), .vss(vss), .out(p[5]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV12_5 ( .in(nbb[5]), .vss(vss), .out(n1[5]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV12_4 ( .in(nbb[4]), .vss(vss), .out(n1[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV12_3 ( .in(nbb[3]), .vss(vss), .out(n1[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV12_2 ( .in(nbb[2]), .vss(vss), .out(n1[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV12_1 ( .in(nbb[1]), .vss(vss), .out(n1[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV12_0 ( .in(nbb[0]), .vss(vss), .out(n1[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV4_3 ( .in(n1[3]), .vss(vss), .out(n[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV4_2 ( .in(n1[2]), .vss(vss), .out(n[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV4_1 ( .in(n1[1]), .vss(vss), .out(n[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV4_0 ( .in(n1[0]), .vss(vss), .out(n[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV6_4 ( .in(p1[4]), .vss(vss), .out(p[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV6_3 ( .in(p1[3]), .vss(vss), .out(p[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV6_2 ( .in(p1[2]), .vss(vss), .out(p[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV6_1 ( .in(p1[1]), .vss(vss), .out(p[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV6_0 ( .in(p1[0]), .vss(vss), .out(p[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV15_5 ( .in(net023[5]), .vss(vss), .out(calp[5]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV15_4 ( .in(net023[4]), .vss(vss), .out(calp[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV15_3 ( .in(net023[3]), .vss(vss), .out(calp[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV15_2 ( .in(net023[2]), .vss(vss), .out(calp[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV15_1 ( .in(net023[1]), .vss(vss), .out(calp[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV15_0 ( .in(net023[0]), .vss(vss), .out(calp[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV16_4 ( .in(net022[4]), .vss(vss), .out(caln[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV16_3 ( .in(net022[3]), .vss(vss), .out(caln[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV16_2 ( .in(net022[2]), .vss(vss), .out(caln[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV16_1 ( .in(net022[1]), .vss(vss), .out(caln[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV16_0 ( .in(net022[0]), .vss(vss), .out(caln[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_SLVT INV14 ( .in(en_up), .vss(vss), .out(enup_b), 
    .vdd(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_6 ( .y(pb[6]), .vss(vss), .vdd(vddq), 
    .b(enup_b), .a(inb_p));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_5 ( .y(pb[5]), .vss(vss), .vdd(vddq), 
    .b(calp[5]), .a(inb_p));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_4 ( .y(pb[4]), .vss(vss), .vdd(vddq), 
    .b(calp[4]), .a(inb_p));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_3 ( .y(pb[3]), .vss(vss), .vdd(vddq), 
    .b(calp[3]), .a(inb_p));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_2 ( .y(pb[2]), .vss(vss), .vdd(vddq), 
    .b(calp[2]), .a(inb_p));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_1 ( .y(pb[1]), .vss(vss), .vdd(vddq), 
    .b(calp[1]), .a(inb_p));

wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt NOR1_0 ( .y(pb[0]), .vss(vss), .vdd(vddq), 
    .b(calp[0]), .a(inb_p));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_7 ( .in(n[5]), .vss(vss), .out(n_fix), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_6 ( .in(n[5]), .vss(vss), .out(n_fix), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_5 ( .in(n[4]), .vss(vss), .out(dn_code[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_4 ( .in(n[4]), .vss(vss), .out(dn_code[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_3 ( .in(n[3]), .vss(vss), .out(dn_code[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_2 ( .in(n[2]), .vss(vss), .out(dn_code[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_1 ( .in(n[1]), .vss(vss), .out(dn_code[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV13_0 ( .in(n[0]), .vss(vss), .out(dn_code[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV17_1 ( .in(n1[5]), .vss(vss), .out(n[5]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV17_0 ( .in(n1[4]), .vss(vss), .out(n[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_8 ( .in(p[6]), .vss(vss), .out(p_fix), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_7 ( .in(p[6]), .vss(vss), .out(p_fix), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_6 ( .in(p[5]), .vss(vss), .out(up_code[5]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_5 ( .in(p[5]), .vss(vss), .out(up_code[5]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_4 ( .in(p[4]), .vss(vss), .out(up_code[4]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_3 ( .in(p[3]), .vss(vss), .out(up_code[3]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_2 ( .in(p[2]), .vss(vss), .out(up_code[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_1 ( .in(p[1]), .vss(vss), .out(up_code[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_SLVT INV9_0 ( .in(p[0]), .vss(vss), .out(up_code[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_240p I8 ( .vddq(vddq), .vss(vss), .out(drv_out), 
    .up_code(up_code), .up_fix(p_fix));

wphy_lp4x5_cmn_NAND2_D1_GL16_SLVT NAND_4 ( .tiehi(vddq), .vdd(vddq), .y(net022[4]), 
    .vss(vss), .tielo(vss), .b(ncal[4]), .a(en_dn));

wphy_lp4x5_cmn_NAND2_D1_GL16_SLVT NAND_3 ( .tiehi(vddq), .vdd(vddq), .y(net022[3]), 
    .vss(vss), .tielo(vss), .b(ncal[3]), .a(en_dn));

wphy_lp4x5_cmn_NAND2_D1_GL16_SLVT NAND_2 ( .tiehi(vddq), .vdd(vddq), .y(net022[2]), 
    .vss(vss), .tielo(vss), .b(ncal[2]), .a(en_dn));

wphy_lp4x5_cmn_NAND2_D1_GL16_SLVT NAND_1 ( .tiehi(vddq), .vdd(vddq), .y(net022[1]), 
    .vss(vss), .tielo(vss), .b(ncal[1]), .a(en_dn));

wphy_lp4x5_cmn_NAND2_D1_GL16_SLVT NAND_0 ( .tiehi(vddq), .vdd(vddq), .y(net022[0]), 
    .vss(vss), .tielo(vss), .b(ncal[0]), .a(en_dn));

wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt NAND0_5 ( .vdd(vddq), .y(nbb[5]), .vss(vss), 
    .b(en_dn), .a(inb_n));

wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt NAND0_4 ( .vdd(vddq), .y(nbb[4]), .vss(vss), 
    .b(caln[4]), .a(inb_n));

wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt NAND0_3 ( .vdd(vddq), .y(nbb[3]), .vss(vss), 
    .b(caln[3]), .a(inb_n));

wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt NAND0_2 ( .vdd(vddq), .y(nbb[2]), .vss(vss), 
    .b(caln[2]), .a(inb_n));

wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt NAND0_1 ( .vdd(vddq), .y(nbb[1]), .vss(vss), 
    .b(caln[1]), .a(inb_n));

wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt NAND0_0 ( .vdd(vddq), .y(nbb[0]), .vss(vss), 
    .b(caln[0]), .a(inb_n));

wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT NOR_5 ( .tiehi(vddq), .tielo(vss), .y(net023[5]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[5]));

wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT NOR_4 ( .tiehi(vddq), .tielo(vss), .y(net023[4]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[4]));

wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT NOR_3 ( .tiehi(vddq), .tielo(vss), .y(net023[3]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[3]));

wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT NOR_2 ( .tiehi(vddq), .tielo(vss), .y(net023[2]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[2]));

wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT NOR_1 ( .tiehi(vddq), .tielo(vss), .y(net023[1]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[1]));

wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT NOR_0 ( .tiehi(vddq), .tielo(vss), .y(net023[0]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[0]));

endmodule
// Library - wphy_gf12lp_lp4x5_sim_lib, Cell - wphy_lp4x5_cmn_tb, View
//- schematic
// LAST TIME SAVED: Jan 17 22:00:01 2021
// NETLIST TIME: Jan 17 22:00:28 2021
`timescale 1ps / 1ps 




 

// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice,
//View - schematic
// LAST TIME SAVED: Dec  2 23:33:43 2020
// NETLIST TIME: Jan 17 22:00:26 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice (out_t, vddq, vss, impd, in_t, ncal, 
    ovrd, ovrd_b, ovrd_n_b, ovrd_p_b, pcal);

output  out_t;

inout  vddq, vss;

input  impd, in_t, ovrd, ovrd_b, ovrd_n_b, ovrd_p_b;

input [4:0]  ncal;
input [5:0]  pcal;


wphy_lp4x5_cmn_wphy_lp4x5_drv_240 I0 ( .pcal(pcal[5:0]), .vddq(vddq), .vss(vss), 
    .drv_out(out_t), .inb_n(data_b), .inb_p(data_b), .ncal(ncal[4:0]), 
    .en_dn(impd), .en_up(impd));

wphy_lp4x5_cmn_wphy_lp4x5_predrv INVT0 ( .pd(ovrd_n_b), .pu(ovrd_p_b), .out(data_b), 
    .en(ovrd_b), .enb(ovrd), .vss(vss), .in(in_t), .vdd(vddq));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_wphy_lp4x5_drv_core, View -
//schematic
// LAST TIME SAVED: Dec 17 15:38:44 2020
// NETLIST TIME: Jan 17 22:00:26 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_wphy_lp4x5_drv_core (out_t, vddq, vss, impd, impd_b, in_t, ncal, 
    ovrd, ovrd_b, ovrd_n_b, ovrd_p_b, pcal);

output  out_t;

inout  vddq, vss;

input  in_t;

input [4:0]  ncal;
input [2:0]  ovrd_p_b;
input [2:0]  ovrd_n_b;
input [2:0]  ovrd_b;
input [2:0]  impd_b;
input [5:0]  pcal;
input [2:0]  ovrd;
input [2:0]  impd;


wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE0 ( .out_t(out_t), .impd(impd[0]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[0]), .ovrd_b(ovrd_b[0]), 
    .ovrd_n_b(ovrd_n_b[0]), .ovrd_p_b(ovrd_p_b[0]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE1_1 ( .out_t(out_t), .impd(impd[1]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[1]), .ovrd_b(ovrd_b[1]), 
    .ovrd_n_b(ovrd_n_b[1]), .ovrd_p_b(ovrd_p_b[1]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE1_0 ( .out_t(out_t), .impd(impd[1]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[1]), .ovrd_b(ovrd_b[1]), 
    .ovrd_n_b(ovrd_n_b[1]), .ovrd_p_b(ovrd_p_b[1]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE2_3 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE2_2 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE2_1 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_core_slice DRV_SLICE2_0 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

endmodule
// Library - wavshared_gf12lp_dig_lib, Cell - wphy_lp4x5_cmn_SE2DIHS_D2_GL16_RVT, View
//- schematic
// LAST TIME SAVED: Jan 12 10:56:44 2021
// NETLIST TIME: Jan 17 22:00:26 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_SE2DIHS_D2_GL16_RVT (outn, outp, vdd, vss, in, tiehi, tielo);

output  outn, outp;

inout  vdd, vss;

input  in, tiehi, tielo;


wphy_lp4x5_cmn_INV_D2_GL16_RVT INV4_1 ( .in(p1), .vss(vss), .out(outn), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV4_0 ( .in(p1), .vss(vss), .out(outn), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV6 ( .in(inb), .vss(vss), .out(p1), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV8 ( .in(in), .vss(vss), .out(inb), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV7 ( .in(in), .vss(vss), .out(inb), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV5_1 ( .in(n1), .vss(vss), .out(outp), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV5_0 ( .in(n1), .vss(vss), .out(outp), .vdd(vdd));

wphy_lp4x5_cmn_PU_D1_GL16_RVT PU0 ( .vdd(vdd), .en(tiehi), .y(inb));

wphy_lp4x5_cmn_PU_D1_GL16_RVT PU1 ( .vdd(vdd), .en(tiehi), .y(n1));

wphy_lp4x5_cmn_XG_D1_GL16_RVT XGATE0_4 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_XG_D1_GL16_RVT XGATE0_3 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_XG_D1_GL16_RVT XGATE0_2 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_XG_D1_GL16_RVT XGATE0_1 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_XG_D1_GL16_RVT XGATE0_0 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_INV_D1_GL16_RVT_Mmod_nomodel INV10 ( .tiehi(tiehi), .tielo(tielo), 
    .in(outp), .vss(vss), .out(outn), .vdd(vdd));

wphy_lp4x5_cmn_INV_D1_GL16_RVT_Mmod_nomodel INV3 ( .tiehi(tiehi), .tielo(tielo), 
    .in(n1), .vss(vss), .out(p1), .vdd(vdd));

wphy_lp4x5_cmn_INV_D1_GL16_RVT_Mmod_nomodel INV2 ( .tiehi(tiehi), .tielo(tielo), 
    .in(p1), .vss(vss), .out(n1), .vdd(vdd));

wphy_lp4x5_cmn_INV_D1_GL16_RVT_Mmod_nomodel INV9 ( .tiehi(tiehi), .tielo(tielo), 
    .in(outn), .vss(vss), .out(outp), .vdd(vdd));

wphy_lp4x5_cmn_PD_D1_GL16_RVT PD0 ( .vss(vss), .enb(tielo), .y(inb));

wphy_lp4x5_cmn_PD_D1_GL16_RVT PD1 ( .vss(vss), .enb(tielo), .y(n1));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_wphy_lp4x5_dq_drvr_w_lpbk,
//View - schematic
// LAST TIME SAVED: Dec 14 16:27:49 2020
// NETLIST TIME: Jan 17 22:00:27 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_wphy_lp4x5_dq_drvr_w_lpbk (d_lpbk_out, rx_in, pad, vdd_aon, 
    vdda, vddq, vss, d_bs_din, d_bs_ena, d_drv_impd, d_in_c, 
    d_lpbk_ena, d_ncal, d_ovrd, d_ovrd_val, d_pcal, freeze_n);

output  d_lpbk_out, rx_in;

inout  pad, vdd_aon, vdda, vddq, vss;

input  d_bs_din, d_bs_ena, d_in_c, d_lpbk_ena, d_ovrd_val, freeze_n;

input [4:0]  d_ncal;
input [5:0]  d_pcal;
input [2:0]  d_ovrd;
input [2:0]  d_drv_impd;

// Buses in the design

wire  [2:0]  impd_b;

wire  [2:0]  ovrd_buf;

wire  [2:0]  net045;

wire  [2:0]  ovrd_b_frz;

wire  [2:0]  impd_b_frz;

wire  [2:0]  ovrd_n_b;

wire  [2:0]  net046;

wire  [2:0]  ovrd_p_b;

wire  [2:0]  ovrd_b;

wire  [2:0]  impd;


wphy_lp4x5_cmn_INV_D8_GL16_RVT INV17_2 ( .in(impd_b[2]), .vss(vss), .out(impd[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D8_GL16_RVT INV17_1 ( .in(impd_b[1]), .vss(vss), .out(impd[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D8_GL16_RVT INV17_0 ( .in(impd_b[0]), .vss(vss), .out(impd[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_drv_core DRV ( .ovrd(ovrd_buf[2:0]), .ovrd_b(ovrd_b[2:0]), 
    .vddq(vddq), .vss(vss), .out_t(pad), .impd(impd[2:0]), 
    .impd_b(impd_b[2:0]), .in_t(in_t), .ncal(d_ncal[4:0]), 
    .ovrd_n_b(ovrd_n_b[2:0]), .ovrd_p_b(ovrd_p_b[2:0]), 
    .pcal(d_pcal[5:0]));

wphy_lp4x5_cmn_wphy_lp4x5_cmn_cdm_50ohm SEC_ESD1 ( .pad(pad), .vdd(vddq), .vss(vss), .out(rx_in));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV16_2 ( .in(impd_b_frz[2]), .vss(vss), 
    .out(net046[2]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV16_1 ( .in(impd_b_frz[1]), .vss(vss), 
    .out(net046[1]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV16_0 ( .in(impd_b_frz[0]), .vss(vss), 
    .out(net046[0]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV15 ( .in(val_b_frz), .vss(vss), .out(net042), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV13_2 ( .in(ovrd_b_frz[2]), .vss(vss), 
    .out(net045[2]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV13_1 ( .in(ovrd_b_frz[1]), .vss(vss), 
    .out(net045[1]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV13_0 ( .in(ovrd_b_frz[0]), .vss(vss), 
    .out(net045[0]), .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV18_2 ( .in(net046[2]), .vss(vss), .out(impd_b[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV18_1 ( .in(net046[1]), .vss(vss), .out(impd_b[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV18_0 ( .in(net046[0]), .vss(vss), .out(impd_b[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV14 ( .in(net042), .vss(vss), .out(ovrd_val_b), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV12_2 ( .in(net045[2]), .vss(vss), .out(ovrd_b[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV12_1 ( .in(net045[1]), .vss(vss), .out(ovrd_b[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV12_0 ( .in(net045[0]), .vss(vss), .out(ovrd_b[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV11_2 ( .in(ovrd_b[2]), .vss(vss), .out(ovrd_buf[2]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV11_1 ( .in(ovrd_b[1]), .vss(vss), .out(ovrd_buf[1]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV11_0 ( .in(ovrd_b[0]), .vss(vss), .out(ovrd_buf[0]), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV10 ( .in(freeze_n), .vss(vss), .out(freeze_vq), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV20 ( .in(bs_enb_vq), .vss(vss), .out(bs_ena_vq), 
    .vdd(vddq));

wphy_lp4x5_cmn_INV_D4_GL16_RVT INV9 ( .in(freeze_vq), .vss(vss), .out(freeze_n_vq), 
    .vdd(vddq));

wphy_lp4x5_cmn_SE2DIHS_D2_GL16_RVT SE2DIFF0 ( .tiehi(vdda), .vdd(vdda), .vss(vss), 
    .tielo(vss), .outp(in_c), .outn(in_t), .in(d_in_c));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND8 ( .tielo(vss), .vdd(vddq), .y(val_b_frz), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd_val));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND3_2 ( .tielo(vss), .vdd(vddq), .y(ovrd_b_frz[2]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd[2]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND3_1 ( .tielo(vss), .vdd(vddq), .y(ovrd_b_frz[1]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd[1]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND0_2 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_b[2]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_val_b), .a(ovrd_buf[2]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND0_1 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_b[1]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_val_b), .a(ovrd_buf[1]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND0_0 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_b[0]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_val_b), .a(ovrd_buf[0]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND4 ( .tielo(vss), .vdd(vddq), .y(bs_data_b), 
    .vss(vss), .tiehi(vddq), .b(freeze_n), .a(d_bs_din));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND5 ( .tielo(vss), .vdd(vddq), .y(bs_enb_vq), 
    .vss(vss), .tiehi(vddq), .b(freeze_n), .a(d_bs_ena));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND1_2 ( .tielo(vss), .vdd(vddq), .y(impd_b_frz[2]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_drv_impd[2]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND1_1 ( .tielo(vss), .vdd(vddq), .y(impd_b_frz[1]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_drv_impd[1]));

wphy_lp4x5_cmn_NOR2_D1_GL16_RVT NOR0_2 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_b[2]), 
    .vss(vss), .vdd(vddq), .b(ovrd_val_b), .a(ovrd_b[2]));

wphy_lp4x5_cmn_NOR2_D1_GL16_RVT NOR0_1 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_b[1]), 
    .vss(vss), .vdd(vddq), .b(ovrd_val_b), .a(ovrd_b[1]));

wphy_lp4x5_cmn_NOR2_D1_GL16_RVT NOR0_0 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_b[0]), 
    .vss(vss), .vdd(vddq), .b(ovrd_val_b), .a(ovrd_b[0]));

wphy_lp4x5_cmn_NOR2_D1_GL16_RVT NAND2 ( .tielo(vss), .tiehi(vddq), .y(impd_b_frz[0]), 
    .vss(vss), .vdd(vddq), .b(freeze_vq), .a(d_drv_impd[0]));

wphy_lp4x5_cmn_NOR2_D1_GL16_RVT NOR1 ( .tielo(vss), .tiehi(vddq), .y(ovrd_b_frz[0]), 
    .vss(vss), .vdd(vddq), .b(freeze_vq), .a(d_ovrd[0]));

wphy_lp4x5_cmn_hbm PRIM_ESD0 ( .vdd(vddq), .vss(vss), .pad(pad));

wphy_lp4x5_cmn_wphy_INVT_D2_GL16_RVT_withR INVT0 ( .out(pad), .en(bs_ena_vq), 
    .enb(bs_enb_vq), .vss(vss), .in(bs_data_b), .vdd(vddq));

wphy_lp4x5_cmn_wphy_lp4x5_lvlsht_vq2va LS0 ( .d_ena(d_lpbk_ena), .vddq(vddq), 
    .out(d_lpbk_out), .outb(net020), .vss(vss), .vdda(vdda), 
    .in_vq(rx_in), .freeze_n(freeze_n));

endmodule
// Library - wavshared_gf12lp_dig_lib, Cell - wphy_lp4x5_cmn_wmx_decoder_3to8_svt,
//View - schematic
// LAST TIME SAVED: Nov 10 12:10:41 2020
// NETLIST TIME: Jan 17 22:00:27 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_wmx_decoder_3to8_svt (y, yb, vdd, vss, a, tiehi, tielo);


inout  vdd, vss;

input  tiehi, tielo;

output [7:0]  yb;
output [7:0]  y;

input [2:0]  a;

// Buses in the design

wire  [2:0]  ab;


wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_7 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[7]), .vss(vss), .c(a[2]), .b(a[1]), .a(a[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_6 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[6]), .vss(vss), .c(a[2]), .b(a[1]), .a(ab[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_5 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[5]), .vss(vss), .c(a[2]), .b(ab[1]), .a(a[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_4 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[4]), .vss(vss), .c(a[2]), .b(ab[1]), .a(ab[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_3 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[3]), .vss(vss), .c(ab[2]), .b(a[1]), .a(a[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_2 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[2]), .vss(vss), .c(ab[2]), .b(a[1]), .a(ab[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_1 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[1]), .vss(vss), .c(ab[2]), .b(ab[1]), .a(a[0]));

wphy_lp4x5_cmn_NAND3_D1_GL16_RVT NAND0_0 ( .tiehi(tiehi), .tielo(tielo), .vdd(vdd), 
    .y(yb[0]), .vss(vss), .c(ab[2]), .b(ab[1]), .a(ab[0]));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_2 ( .in(a[2]), .vss(vss), .out(ab[2]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_1 ( .in(a[1]), .vss(vss), .out(ab[1]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_0 ( .in(a[0]), .vss(vss), .out(ab[0]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_7 ( .in(yb[7]), .vss(vss), .out(y[7]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_6 ( .in(yb[6]), .vss(vss), .out(y[6]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_5 ( .in(yb[5]), .vss(vss), .out(y[5]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_4 ( .in(yb[4]), .vss(vss), .out(y[4]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_3 ( .in(yb[3]), .vss(vss), .out(y[3]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_2 ( .in(yb[2]), .vss(vss), .out(y[2]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_1 ( .in(yb[1]), .vss(vss), .out(y[1]), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV_0 ( .in(yb[0]), .vss(vss), .out(y[0]), .vdd(vdd));

endmodule
// Library - wavshared_gf12lp_dig_lib, Cell - wphy_lp4x5_cmn_MUXATEST_D2_GL150_EG,
//View - schematic
// LAST TIME SAVED: Nov 24 10:17:09 2020
// NETLIST TIME: Jan 17 22:00:27 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_MUXATEST_D2_GL150_EG (atst_out, vdd, vdda1p8, vss, freezeb_hv, 
    in, sel);

output  atst_out;

inout  vdd, vdda1p8, vss;

input  freezeb_hv;

input [7:1]  in;
input [2:0]  sel;

// Buses in the design

wire  [7:0]  selhb;

wire  [7:0]  selh;

wire  [7:0]  s;

wire  [7:0]  net4;


wphy_lp4x5_cmn_wmx_decoder_3to8_svt DECODER3to8 ( .vdd(vdd), .y(s[7:0]), 
    .yb(net4[7:0]), .a(sel[2:0]), .tielo(tielo), .tiehi(tiehi), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_7 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[7]), .in(s[7]), .outp(selh[7]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_6 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[6]), .in(s[6]), .outp(selh[6]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_5 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[5]), .in(s[5]), .outp(selh[5]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_4 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[4]), .in(s[4]), .outp(selh[4]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_3 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[3]), .in(s[3]), .outp(selh[3]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_2 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[2]), .in(s[2]), .outp(selh[2]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_1 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[1]), .in(s[1]), .outp(selh[1]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0_0 ( .freezeb_hv(freezeb_hv), 
    .outn(selhb[0]), .in(s[0]), .outp(selh[0]), .vdda1p8(vdda1p8), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_0 ( .vdda1p8(vdda1p8), .out(atst_out), 
    .en(selhb[0]), .enb(selh[0]), .in(o1), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_7 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[7]), 
    .enb(selhb[7]), .in(in[7]), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_6 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[6]), 
    .enb(selhb[6]), .in(in[6]), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_5 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[5]), 
    .enb(selhb[5]), .in(in[5]), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_4 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[4]), 
    .enb(selhb[4]), .in(in[4]), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_3 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[3]), 
    .enb(selhb[3]), .in(in[3]), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_2 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[2]), 
    .enb(selhb[2]), .in(in[2]), .vss(vss));

wphy_lp4x5_cmn_XG_D2_GL150_EG XG0_1 ( .vdda1p8(vdda1p8), .out(o1), .en(selh[1]), 
    .enb(selhb[1]), .in(in[1]), .vss(vss));

wphy_lp4x5_cmn_TIELO_D2_GL16_RVT I2 ( .tielo(tielo), .vss(vss), .vdd(vdd));

wphy_lp4x5_cmn_TIEHI_D2_GL16_RVT I3 ( .tiehi(tiehi), .vss(vss), .vdd(vdd));

endmodule
// Library - wavshared_gf12lp_dig_lib, Cell -
//wphy_lp4x5_cmn_MUXATEST_D2_14to1_GL150_EG, View - schematic
// LAST TIME SAVED: Nov 10 11:37:44 2020
// NETLIST TIME: Jan 17 22:00:27 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_MUXATEST_D2_14to1_GL150_EG (atst_out, vdd, vdda1p8, vss, 
    atst_sel, freezeb_hv, in);

output  atst_out;

inout  vdd, vdda1p8, vss;

input  freezeb_hv;

input [3:0]  atst_sel;
input [13:0]  in;

// Buses in the design

wire  [2:0]  sel0;

wire  [2:0]  net47;

wire  [2:0]  net46;

wire  [2:0]  sel1;


wphy_lp4x5_cmn_MUXATEST_D2_GL150_EG ATST0 ( .vdda1p8(vdda1p8), 
    .freezeb_hv(freezeb_hv), .atst_out(atst_out), .in(in[6:0]), 
    .sel(sel0[2:0]), .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_MUXATEST_D2_GL150_EG ATST1 ( .vdda1p8(vdda1p8), 
    .freezeb_hv(freezeb_hv), .atst_out(atst_out), .in(in[13:7]), 
    .sel(sel1[2:0]), .vdd(vdd), .vss(vss));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND1_2 ( .tielo(tielo), .vdd(vdd), .y(net46[2]), 
    .vss(vss), .tiehi(tiehi), .b(sel3b), .a(atst_sel[2]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND1_1 ( .tielo(tielo), .vdd(vdd), .y(net46[1]), 
    .vss(vss), .tiehi(tiehi), .b(sel3b), .a(atst_sel[1]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND1_0 ( .tielo(tielo), .vdd(vdd), .y(net46[0]), 
    .vss(vss), .tiehi(tiehi), .b(sel3b), .a(atst_sel[0]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND0_2 ( .tielo(tielo), .vdd(vdd), .y(net47[2]), 
    .vss(vss), .tiehi(tiehi), .b(atst_sel[3]), .a(atst_sel[2]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND0_1 ( .tielo(tielo), .vdd(vdd), .y(net47[1]), 
    .vss(vss), .tiehi(tiehi), .b(atst_sel[3]), .a(atst_sel[1]));

wphy_lp4x5_cmn_NAND2_D1_GL16_RVT NAND0_0 ( .tielo(tielo), .vdd(vdd), .y(net47[0]), 
    .vss(vss), .tiehi(tiehi), .b(atst_sel[3]), .a(atst_sel[0]));

wphy_lp4x5_cmn_TIEHI_D2_GL16_RVT I0 ( .tiehi(tiehi), .vss(vss), .vdd(vdd));

wphy_lp4x5_cmn_TIELO_D2_GL16_RVT I1 ( .tielo(tielo), .vss(vss), .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV2 ( .in(atst_sel[3]), .vss(vss), .out(sel3b), 
    .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_2 ( .in(net47[2]), .vss(vss), .out(sel1[2]), 
    .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_1 ( .in(net47[1]), .vss(vss), .out(sel1[1]), 
    .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_0 ( .in(net47[0]), .vss(vss), .out(sel1[0]), 
    .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_2 ( .in(net46[2]), .vss(vss), .out(sel0[2]), 
    .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_1 ( .in(net46[1]), .vss(vss), .out(sel0[1]), 
    .vdd(vdd));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_0 ( .in(net46[0]), .vss(vss), .out(sel0[0]), 
    .vdd(vdd));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn, View -
//schematic
// LAST TIME SAVED: Jan 14 14:43:54 2021
// NETLIST TIME: Jan 17 22:00:28 2021
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_lp4x5_cmn (ddr_rstn_lpbk_out, freeze_n_aon, freeze_n_hv, 
    pmon_nand_fout, pmon_nor_fout, vref, zacal_comp_out, pad_atb, 
    pad_reset_n, pad_rext,      
    atst_in, atst_sel, ddr_rstn_bs_din, ddr_rstn_bs_ena, ddr_rstn_din, 
    ddr_rstn_lpbk_ena, dtst_drv_impd, dtst_in, freeze_n, ldo_atst_sel, 
    ldo_phy_ena, ldo_phy_hiz, ldo_tran_enh_ena, ldo_vref_ctrl, 
    pmon_nand_ena, pmon_nor_ena, vref_ctrl, vref_ena, vref_hiz, 
    vref_pwr, zqcal_cal_ena, zqcal_ncal, zqcal_pcal, zqcal_pd_sel, 
    zqcal_vol_0p6_sel
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda1p2  
 ,vddq  
 ,vdd_phy  
 ,vdd_aon  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda1p2;
assign vdda1p2=1'b1;
wire vddq;
assign vddq=1'b1;
wire vdd_phy;
assign vdd_phy=1'b1;
wire vdd_aon;
assign vdd_aon=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda1p2;
inout vddq;
inout vdd_phy;
inout vdd_aon;
inout vss;
`endif


output  ddr_rstn_lpbk_out, freeze_n_aon, freeze_n_hv, pmon_nand_fout, 
    pmon_nor_fout, vref, zacal_comp_out;

inout  pad_atb, pad_reset_n, pad_rext;

input  ddr_rstn_bs_din, ddr_rstn_bs_ena, ddr_rstn_din, 
    ddr_rstn_lpbk_ena, dtst_in, freeze_n, ldo_phy_ena, ldo_phy_hiz, 
    ldo_tran_enh_ena, pmon_nand_ena, pmon_nor_ena, vref_ena, vref_hiz, 
    zqcal_cal_ena, zqcal_pd_sel, zqcal_vol_0p6_sel;

input [2:0]  dtst_drv_impd;
input [1:0]  vref_pwr;
input [5:0]  zqcal_pcal;
input [7:0]  vref_ctrl;
input [4:0]  zqcal_ncal;
input [7:0]  ldo_vref_ctrl;
input [2:0]  ldo_atst_sel;
input [3:0]  atst_in;
input [3:0]  atst_sel;

// Buses in the design 
`ifdef SYNTHESIS 
`else

wire  [7:0]  net1;

wire  [1:0]  net0165;

wire  [1:0]  net0169;

wire  [5:0]  net0168;

wire  [7:0]  vref_ctrl_hv;

wire  [2:0]  ldo_atst_sel_hv;

wire  [7:0]  ldo_ref_ctrl_hv;

wire  [2:0]  net0167;

wire  [1:0]  vref_pwr_hv;


wphy_lp4x5_cmn_wphy_lp4x5_refgen_hv_v3 REFGEN ( .vref_ctrl_hv(vref_ctrl_hv), 
    .vddq(vddq), .vref(vref), .hiz_hv(vref_hiz_hv), 
    .pwr_hv(vref_pwr_hv), .ena_hv(vref_ena_hv), .vss(vss), 
    .vdda1p2(vdda1p2));

wphy_lp4x5_cmn_wphy_lp4x5_zq_cal ZQCAL ( .pad_rext(pad_rext), .vdda(vdd_aon), 
    .vddq(vddq), .vss(vss), .d_cal_comp_out(zacal_comp_out), 
    .d_cal_ena(zqcal_cal_ena), .d_ncal(zqcal_ncal), 
    .d_pcal(zqcal_pcal), .d_pd_sel(zqcal_pd_sel), 
    .d_voh_0p6_sel(zqcal_vol_0p6_sel));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_7 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_6 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_5 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_4 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_3 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_2 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_1 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_INV_D1_GL150_EGU INV2_0 ( .vdda1p2(vdda1p2), .in(net0150), .vss(vss), 
    .out(freeze_n_hv));

wphy_lp4x5_cmn_wphy_pmon_svt_nand PMON_NAND ( .pmon_fout(pmon_nand_fout), 
    .vdda(vdd_phy), .vss(vss), .pmon_en(pmon_nand_ena));

wphy_lp4x5_cmn_LVLHC1_D1_GL16_RVT LVLSFT9_1 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0169[1]), .in(ldo_vref_ctrl[6]), 
    .outp(ldo_ref_ctrl_hv[6]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC1_D1_GL16_RVT LVLSFT9_0 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0169[0]), .in(ldo_vref_ctrl[4]), 
    .outp(ldo_ref_ctrl_hv[4]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_wphy_lp4x5_cke_drvr_w_lpbk IRST_N_DRV ( .d_in_c(ddr_rstn_din), 
    .d_bs_din(ddr_rstn_bs_din), .d_bs_ena(ddr_rstn_bs_ena), 
    .freeze_n_hv(freeze_n_hv), .d_lpbk_out(ddr_rstn_lpbk_out), 
    .pad_cke_out(pad_reset_n), .d_lpbk_ena(ddr_rstn_lpbk_ena), 
    .d_ovrd({vss, vss, vss}), .d_ovrd_val(vss), .vdda(vdd_aon), 
    .vdda1p2(vdda1p2), .vss(vss));

wphy_lp4x5_cmn_wphy_lp4x5_dq_drvr_w_lpbk DTST_DRV ( .vdd_aon(vdd_aon), .d_bs_ena(vss), 
    .rx_in(atest), .d_in_c(dtst_in), .d_lpbk_ena(vss), 
    .freeze_n(freeze_n), .d_lpbk_out(d_lpbk_out), .vdda(vdd_aon), 
    .vddq(vddq), .vss(vss), .d_bs_din(vss), 
    .d_drv_impd(dtst_drv_impd[2:0]), .pad(pad_atb), 
    .d_ncal(zqcal_ncal[4:0]), .d_ovrd({vss, vss, vss}), 
    .d_ovrd_val(vss), .d_pcal(zqcal_pcal[5:0]));

wphy_lp4x5_cmn_wphy_pmon_svt_nor PMON_NOR ( .vdda(vdd_phy), .vss(vss), 
    .pmon_fout(pmon_nor_fout), .pmon_en(pmon_nor_ena));

wire ldo_atst_out_hv;

wphy_lp4x5_cmn_MUXATEST_D2_14to1_GL150_EG GLBL_ATST ( .atst_out(atest), 
    .atst_sel(atst_sel[3:0]), .freezeb_hv(freeze_n_int_hv), 
    .in({atst_in[3:0], ldo_atst_out_hv, vss, vss, vss, vss, vss, vss, 
    vss, vss, vss}), .vss(vss), .vdda1p8(vdda1p2), .vdd(vdd_aon));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT10 ( .freezeb_hv(vdda1p2), .outn(net0150), 
    .in(freeze_n_aon), .outp(freeze_n_int_hv), .vdda1p8(vdda1p2), 
    .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT2_5 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0168[5]), .in(ldo_vref_ctrl[7]), 
    .outp(ldo_ref_ctrl_hv[7]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT2_4 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0168[4]), .in(ldo_vref_ctrl[5]), 
    .outp(ldo_ref_ctrl_hv[5]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT2_3 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0168[3]), .in(ldo_vref_ctrl[3]), 
    .outp(ldo_ref_ctrl_hv[3]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT2_2 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0168[2]), .in(ldo_vref_ctrl[2]), 
    .outp(ldo_ref_ctrl_hv[2]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT2_1 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0168[1]), .in(ldo_vref_ctrl[1]), 
    .outp(ldo_ref_ctrl_hv[1]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT2_0 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0168[0]), .in(ldo_vref_ctrl[0]), 
    .outp(ldo_ref_ctrl_hv[0]), .vdda1p8(vdda1p2), .vdd(vdd_aon), 
    .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT0 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0153), .in(ldo_tran_enh_ena), .outp(ldo_tran_enh_ena_hv), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT4 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0156), .in(ldo_phy_ena), .outp(phy_ena_hv), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT8_2 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0167[2]), .in(ldo_atst_sel[2]), .outp(ldo_atst_sel_hv[2]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT8_1 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0167[1]), .in(ldo_atst_sel[1]), .outp(ldo_atst_sel_hv[1]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT8_0 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0167[0]), .in(ldo_atst_sel[0]), .outp(ldo_atst_sel_hv[0]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT6 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0155), .in(ldo_phy_hiz), .outp(phy_hiz_hv), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT7_1 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0165[1]), .in(vref_pwr[1]), .outp(vref_pwr_hv[1]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT7_0 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0165[0]), .in(vref_pwr[0]), .outp(vref_pwr_hv[0]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT3 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0158), .in(vref_ena), .outp(vref_ena_hv), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_7 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[7]), .in(vref_ctrl[7]), .outp(vref_ctrl_hv[7]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_6 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[6]), .in(vref_ctrl[6]), .outp(vref_ctrl_hv[6]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_5 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[5]), .in(vref_ctrl[5]), .outp(vref_ctrl_hv[5]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_4 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[4]), .in(vref_ctrl[4]), .outp(vref_ctrl_hv[4]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_3 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[3]), .in(vref_ctrl[3]), .outp(vref_ctrl_hv[3]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_2 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[2]), .in(vref_ctrl[2]), .outp(vref_ctrl_hv[2]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_1 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[1]), .in(vref_ctrl[1]), .outp(vref_ctrl_hv[1]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT5_0 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net1[0]), .in(vref_ctrl[0]), .outp(vref_ctrl_hv[0]), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT LVLSFT1 ( .freezeb_hv(freeze_n_int_hv), 
    .outn(net0157), .in(vref_hiz), .outp(vref_hiz_hv), 
    .vdda1p8(vdda1p2), .vdd(vdd_aon), .vss(vss));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_3 ( .in(freeze_n), .vss(vss), .out(freeze_nb), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_2 ( .in(freeze_n), .vss(vss), .out(freeze_nb), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_1 ( .in(freeze_n), .vss(vss), .out(freeze_nb), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV0_0 ( .in(freeze_n), .vss(vss), .out(freeze_nb), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_7 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_6 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_5 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_4 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_3 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_2 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_1 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

wphy_lp4x5_cmn_INV_D2_GL16_RVT INV1_0 ( .in(freeze_nb), .vss(vss), .out(freeze_n_aon), 
    .vdd(vdd_aon));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else



 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_TIEHI_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_TIEHI_D2_GL16_RVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);


  output tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tiehi = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tiehi =  1'b1 ;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_TIELO_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_TIELO_D2_GL16_RVT ( tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  output tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tielo = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tielo =  1'b0 ;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "XG_D2_GL150_18" "systemVerilog"


module wphy_lp4x5_cmn_XG_D2_GL150_EG ( out, en, enb, in
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdda1p8 
`endif //WLOGIC_MODEL_NO_PG
); 

  input in;
  output out;
  input en;
  input enb;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p8;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdda1p8;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

assign out = (en && ~enb) ? in:1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_NAND3_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_NAND3_D1_GL16_RVT ( y, a, b, c
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input c;
  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b&c);

endmodule
//Verilog HDL for "wmx_prs_lib", "wmx_prs_pmon_lvt" "functional"

`timescale 1ns/1ps
module wphy_lp4x5_cmn_wphy_pmon_svt_nor ( pmon_fout, vdda, vss, pmon_en );

  inout vdda;
  input pmon_en;
  output pmon_fout;
  inout vss;

  wire pg_en;
  assign pg_en = vdda & ~vss  ;

  reg fout_pre;
  real PMON_DELAY =1.428571; //in ns, 1.25 for 800MHZ
  real ldo_out_real = 800.0;

initial begin

`ifdef WPHY_LDO_MODEL_INCLUDED
   ldo_out_real = ILDO_PHY.VREFGEN.vref_mv*1e-3;
`else
   ldo_out_real = 800.0*1e-3;
`endif
   PMON_DELAY =  (8.53445*ldo_out_real*ldo_out_real - 16.821*ldo_out_real+9.3735);
   fout_pre = 1'b0;
   #10 fout_pre = 1'b1;
end

always @(posedge fout_pre) begin
`ifdef WPHY_LDO_MODEL_INCLUDED
   ldo_out_real = ILDO_PHY.VREFGEN.vref_mv*1e-3;
`else
   ldo_out_real = 800.0*1e-3;
`endif
   PMON_DELAY =   (8.53445*ldo_out_real*ldo_out_real - 16.821*ldo_out_real+9.3735);
   #(0.5*PMON_DELAY) fout_pre <= ~fout_pre;
   #(0.5*PMON_DELAY) fout_pre <= ~fout_pre;
end

assign pmon_fout = pg_en ? (fout_pre & pmon_en) : 1'bx; 

endmodule
//Verilog HDL for "wphy_lp4x5_lib", "wphy_lp4x5_cmn_wphy_lp4x5_lvlsht_vq2va" "functional"


module wphy_lp4x5_cmn_wphy_lp4x5_lvlsht_vq2va ( out, outb, vdda, vddq, vss, d_ena, freeze_n, in_vq );

  inout vdda;
  output out;
  input in_vq;
  input d_ena;
  input freeze_n;
  output outb;
  inout vddq;
  inout vss;

  wire out_int;

  wire check_en;

`ifdef WANALOG_CHECK_VALID_OUT
  assign check_en=1'b1;
`else
  assign check_en=1'b0;
`endif

	wire pwr_ok;
	assign pwr_ok = vdda & freeze_n &vddq & ~vss;
   assign out_int = pwr_ok ? (in_vq &d_ena ):1'bx;
   assign out  = (check_en===1'b1 && out_int===1'bx) ? 1'b1 : out_int;    // FIXME: ADDED per Sushma's request, may remove it later
	assign outb = ~out;

//   wire pwr_ok;
//   assign pwr_ok = vdda & freeze_n &vddq & ~vss;
//   assign out = pwr_ok ? (in_vq &d_ena ):1'bx;
//   assign outb = ~out;
endmodule
//Verilog HDL for "Serdes", "cmos_inv2_tst" "behavioral"


module wphy_lp4x5_cmn_wphy_INVT_D2_GL16_RVT_withR( in, vdd, vss, out, en, enb );

  inout vss;
  input in;
  inout vdd;
  input en, enb;
  output out;
  wire out;

assign out= (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule



module wphy_lp4x5_cmn_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_PD_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_cmn_PD_D1_GL16_RVT( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_INV_D1_GL16_RVT_Mmod_nomodel"
//"systemVerilog"


module wphy_lp4x5_cmn_INV_D1_GL16_RVT_Mmod_nomodel ( in, out, tiehi, tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
  input tiehi;
  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_XG_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_XG_D1_GL16_RVT ( y, en, enb, a
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input a;
  input en;
  output y;
  input enb;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign y = (en && ~enb) ? a:1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_PU_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_PU_D1_GL16_RVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_INV_D4_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_INV_D4_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;


endmodule
//systemVerilog HDL for "wavshared_gf12lp_ana_lib", "wphy_lp4x5_cmn_cdm" "systemVerilog"

module wphy_lp4x5_cmn_wphy_lp4x5_cmn_cdm_50ohm ( out, pad, vdd, vss );

  inout pad;
  inout vdd;
  inout out;
  inout vss;


wire power_ok;
assign power_ok = vdd & (~vss);

assign pad = power_ok ? out : 1'bx;

endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_cmn_wphy_lp4x5_predrv" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_cmn_wphy_lp4x5_predrv ( out, vdd, vss, en, enb, in, pd, pu );

  input in;
  input pu;
  output out;
  input en;
  inout vdd;
  input pd;
  input enb;
  inout vss;

wire power_ok;
assign power_ok = ~vss & vdd;

assign #(10) out= power_ok ? (en) ? ~in:1'bz : 1'bx;
assign #(10) out= (pu) ? 1'bz:1'b1;
assign #(10) out= (pd) ? 1'b0:1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_NOR2_D1_GL16_SLVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//Verilog HDL for "wavshared_tsmc14lpp_lib", "wphy_lp4x5_cmn_NAND2_D1_GL16_RVT" "functional"


module wphy_lp4x5_cmn_wphy_lp4x5_nanad_d2_slvt ( y, a, b, vdd, vss );

  input b;
  input a;
  inout vdd;
  output y;
  inout vss;


assign y=~(a&b);


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "NAND2_D1_GL16_LVT" "systemVerilog"


module wphy_lp4x5_cmn_NAND2_D1_GL16_SLVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//Verilog HDL for "wmx_lpddr5_lib", "wmx_lpddr5_drv_240p" "functional"


module wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_240p ( out, vddq, vss, up_code, up_fix );

  input up_fix;
  output out;
  inout vddq;
  input  [5:0] up_code;
  inout vss;

  wire power_ok;
  assign power_ok = vddq & ~vss ;
  wire in_ok;
  assign in_ok = (up_code <63) == (~up_fix);
  wire  inb_pn ;
  assign inb_pn = (power_ok&in_ok) ?  ~up_fix   : 1'bx;
  

  assign (supply1, weak0) out = 	(inb_pn == 1'b1 ) ? 1'b1: 	
						 		(inb_pn == 1'b0 ) ? 1'bz : 1'bx ;
endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_INV_D4_GL16_SLVT" "systemVerilog"


module wphy_lp4x5_cmn_INV_D4_GL16_SLVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;


endmodule
//Verilog HDL for "wavshared_tsmc14lpp_lib", "wphy_lp4x5_cmn_NOR2_D1_GL16_RVT" "functional"


module wphy_lp4x5_cmn_wphy_lp4x5_nor_d2_slvt ( y, a, b, vdd, vss );

  input b;
  input a;
  inout vdd;
  output y;
  inout vss;

assign y=~(a|b);
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "INV_D2_GL16_LVT" "systemVerilog"

module wphy_lp4x5_cmn_INV_D2_GL16_SLVT( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_INV_D1_GL16_SLVT" "systemVerilog"

module wphy_lp4x5_cmn_INV_D1_GL16_SLVT( in, out
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign out = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out =  ~in;

endmodule
//Verilog HDL for "wmx_lpddr5_lib", "wmx_lpddr5_drv_240n" "functional"


module wphy_lp4x5_cmn_wphy_lp4x5_cmn_wphy_lp4x5_drv_240n ( out, dn_code, dn_fix, vss );

  input dn_fix;
  output out;
  input  [4:0] dn_code;
  inout vss;


  wire power_ok;
  assign power_ok =  ~vss ;
  wire in_ok;
  assign in_ok = (dn_code >0) == (dn_fix);
  wire  inb_pn ;
  assign inb_pn = (power_ok&in_ok) ?  dn_fix   : 1'bx;
  

  assign (supply1, weak0) out = 	(inb_pn == 1'b1 ) ? 1'b0: 	
						 		(inb_pn == 1'b0 ) ? 1'bz : 1'bx ;


endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_INV_D8_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_INV_D8_GL16_RVT ( in,  out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "NAND2_D1_GL150_UD12" "systemVerilog"


module wphy_lp4x5_cmn_NAND2_D1_GL150_EGU ( y, a, b
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdda1p2 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p2;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdda1p2;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y = ~(a&b);


endmodule
//Verilog HDL for "wavshared_gf12lp_ana_lib", "wphy_lp4x5_cmn_hbm" "functional"


module wphy_lp4x5_cmn_hbm ( pad, vdd, vss );

  inout pad;
  inout vdd;
  inout vss;
endmodule
//systemVerilog HDL for "wavshared_gf12lp_ana_lib", "wphy_lp4x5_cmn_cdm" "systemVerilog"
`timescale 1ps/1ps
module wphy_lp4x5_cmn_cdm ( out, pad, vdd, vss );

  inout out;
  inout vdd;
  inout pad;
  inout vss;

string str_out;
string str_pad;
reg assert_en=1'b0;

wire power_ok;
assign power_ok = vdd & (~vss);
assign (weak1, weak0) pad = power_ok ? out : 1'bx;
assign (weak1, weak0) out = power_ok ? pad : 1'bx;

initial begin
   if ($value$plusargs("WPHY_ANA_ASSERT_EN=%f", assert_en)) begin
      assert_en=assert_en;
   end
end


always @(out,pad) begin
   if(assert_en) begin
      str_out = $sformatf("%v", out);
      //$display("out strength=%s",str_out);
      str_pad = $sformatf("%v", pad);
      //$display("pad strength=%s",str_pad);

      if(((str_pad=="St1") || (str_pad=="St0")) && ((str_out=="St0") || (str_out=="St1"))) begin
         $display(" WPHY_ANA_ERROR: potential contention, ports driven from both sides in %m at %t",$realtime);
      end
   end
end

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_NOR3_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_NOR3_D1_GL16_RVT ( y, a, b, c
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input c;
  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y = ~(a|b|c);



endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_LVLHC0_D1_GL16_RVT ( outn, outp, in, freezeb_hv
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd, vdda1p8 
`endif //WLOGIC_MODEL_NO_PG
); 

  input freezeb_hv;
  input in;
  output outn;
  output outp;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p8;
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
  assign outp = ~freezeb_hv ? 1'b0 : in;
  assign outn = ~freezeb_hv ? 1'b1 : ~in;
`else

  assign outp = (vdd & vdda1p8 & ~vss) ? (~freezeb_hv ? 1'b0 : in)  : 1'b0;
  assign outn = (vdd & vdda1p8 & ~vss) ? (~freezeb_hv ? 1'b1 : ~in) : 1'b0;

`endif //WLOGIC_MODEL_NO_PG



endmodule
//Verilog HDL for "wphy_lp4x5_lib", "wphy_lp4x5_cmn_wphy_lp4x5_cke_drv_core" "functional"


module wphy_lp4x5_cmn_wphy_lp4x5_cke_drv_core ( out_h, vdda1p2, vss, inb_h );

  output out_h;
  inout vdda1p2;
  input inb_h;
  inout vss;

	wire pwr_ok;
	assign pwr_ok = vdda1p2 & ~vss;
	assign out_h = pwr_ok ? ~inb_h : 1'bx;
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_NOR2_D1_GL16_LVT" "systemVerilog"


module wphy_lp4x5_cmn_NOR2_D1_GL16_LVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_INV_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_MUXT2_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_MUXT2_D2_GL16_RVT( yb, a, b, s, sb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input a; 
  input sb;
  input s;
  output yb;
  input b;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire yb;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign yb = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign yb = (s && ~sb) ? ~b:~a;



endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_LVLHC1_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_LVLHC1_D1_GL16_RVT ( outn, outp, in, freezeb_hv
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd, vdda1p8 
`endif //WLOGIC_MODEL_NO_PG
); 

  input freezeb_hv;
  input in;
  output outn;
  output outp;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p8;
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
  assign outp = ~freezeb_hv ? 1'b0 : in;
  assign outn = ~freezeb_hv ? 1'b1 : ~in;
`else

  assign outp = (vdd & vdda1p8 & ~vss) ? (~freezeb_hv ? 1'b1 : in)  : 1'b0;
  assign outn = (vdd & vdda1p8 & ~vss) ? (~freezeb_hv ? 1'b0 : ~in) : 1'b0;

`endif //WLOGIC_MODEL_NO_PG



endmodule
//Verilog HDL for "wmx_prs_lib", "wmx_prs_pmon_lvt" "functional"

`timescale 1ns/1ps
module wphy_lp4x5_cmn_wphy_pmon_svt_nand ( pmon_fout, vdda, vss, pmon_en );

  inout vdda;
  input pmon_en;
  output pmon_fout;
  inout vss;

  wire pg_ok;
  assign pg_ok = vdda & ~vss ;

  reg fout_pre;
  real PMON_DELAY = 1.42857; //in ns, 1.25 for 800MHZ
  real ldo_out_real = 800.0;  //800mV

initial begin

`ifdef WPHY_LDO_MODEL_INCLUDED
   ldo_out_real = ILDO_PHY.VREFGEN.vref_mv*1e-3;
`else
   ldo_out_real = 800.0*1e-3;
`endif
   PMON_DELAY =  (7.8585*ldo_out_real*ldo_out_real - 15.636*ldo_out_real+8.9138);
   fout_pre = 1'b0;
   #10 fout_pre = 1'b1;
end

always @(posedge fout_pre) begin
`ifdef WPHY_LDO_MODEL_INCLUDED
   ldo_out_real = ILDO_PHY.VREFGEN.vref_mv*1e-3;
`else
   ldo_out_real = 800.0*1e-3;
`endif
   PMON_DELAY =  (7.8585*ldo_out_real*ldo_out_real - 15.636*ldo_out_real+8.9138);
   #(0.5*PMON_DELAY) fout_pre <= ~fout_pre;
   #(0.5*PMON_DELAY) fout_pre <= ~fout_pre;
end

assign pmon_fout = pg_ok ? (fout_pre & pmon_en) : 1'bx; 

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "INV_D1_GL150_UD12" "systemVerilog"


module wphy_lp4x5_cmn_INV_D1_GL150_EGU ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdda1p2, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p2;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdda1p2;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wmx_lpddr5_lib", "wmx_lpddr5_ZQ_cal" "systemVerilog"


module wphy_lp4x5_cmn_wphy_lp4x5_zq_cal ( d_cal_comp_out, pad_rext, vdda, vddq, vss, d_cal_ena,
d_ncal, d_pcal, d_pd_sel, d_voh_0p6_sel );

  input d_pd_sel;
  input d_voh_0p6_sel;
  input d_cal_ena;
  inout vdda;
 // input ip25u_n;
  input  [4:0] d_ncal;
  inout vddq;
  inout pad_rext;
  output reg d_cal_comp_out;
  input  [5:0] d_pcal;
  inout vss;

real Rfix_n = 500;
real Rfix_p =  1000;
real Rn = 7400;
real Rp = 6000;
real vq =0.5;
real Vq_mV;
real Rpd, Rpu, Vpd, Vpu, vin, vref;
wire pwr_ok;

assign pwr_ok = (~vss &vdda &vddq);

initial begin

	if ($value$plusargs("VDDQ=%f",Vq_mV)) begin
		vq = Vq_mV/1000; 
	end else begin 
		vq = 0.5;
	end
	Rpd = 1/(1/Rfix_n +d_ncal/Rn);
	Rpu = 1/(1/Rfix_p +~d_pcal/Rp);
	Vpd = vq*Rpd/(240+Rpd);
	Vpu = vq*Rpd/(Rpd+Rpu);
	vref = d_pd_sel? 0.5*vq : (d_voh_0p6_sel? 0.6*vq : 0.5*vq);
	vin  = d_pd_sel ? Vpd : Vpu;
	d_cal_comp_out =  pwr_ok ? (~d_cal_ena ? 1'b0 : (vin > vref ? 1'b1 : 1'b0)):1'bx;
end
always @(d_pcal or d_ncal or d_cal_ena or d_pd_sel or d_voh_0p6_sel ) begin
	Rpd = 1/(1/Rfix_n +d_ncal/Rn);
	Rpu = 1/(1/Rfix_p +~d_pcal/Rp);
	Vpd = vq*Rpd/(240+Rpd);
	Vpu = vq*Rpd/(Rpd+Rpu);
	vref = d_pd_sel? 0.5*vq : (d_voh_0p6_sel? 0.6*vq : 0.5*vq);
	vin  = d_pd_sel ? Vpd : Vpu;
	d_cal_comp_out =  pwr_ok ? (~d_cal_ena ? 1'b0 : (vin > vref ? 1'b1 : 1'b0)):1'bx;
end
endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_cmn_wphy_lp4x5_refgen_hv_v3" "systemVerilog"

`timescale 1ns/1ps

module wphy_lp4x5_cmn_wphy_lp4x5_refgen_hv_v3 ( vref, vdda1p2, vddq, vss, ena_hv, hiz_hv, pwr_hv,
vref_ctrl_hv );

  input ena_hv;
  input  [7:0] vref_ctrl_hv;
`ifdef WPIN_EN
  output integer vref;
`else
  output vref;
`endif
  input  [1:0] pwr_hv;
  inout vddq;
  inout vdda1p2;
  input hiz_hv;
  inout vss;

`ifdef WPIN_EN
`elsif WPIN_UART_EN
Wpin_uart_tx Wvref(vref);
`else
  reg vref=1'b0;
`endif

wire pwr_ok;
var integer b2d_v =0;
var  integer val ; //in mv
integer i ;
//integer step = 2;//2mv
integer offset = 0;//50mv offset 

real dly_ns = 10; //in ns
integer step =2 ; //in mv

assign pwr_ok= ~vss & vdda1p2 & vddq;
initial begin
   dly_ns = pwr_hv*10 +10;
end

always @(*) begin
   dly_ns = pwr_hv*10 +10;
   val = vref_ctrl_hv*step+offset;
   if (pwr_ok) begin
      if (hiz_hv) begin
`ifdef WPIN_UART_EN
         Wvref.en=1'b0;
`else
         vref= 1'bZ;
`endif   
      end else if (ena_hv) begin
`ifdef WPIN_EN
         #dly_ns vref = val;
`elsif WPIN_UART_EN
         Wvref.en=1'b1;
         #dly_ns;
         Wvref.value=val;
`else
         #dly_ns vref = 1'b1;
`endif
      end 
      else begin
`ifdef WPIN_UART_EN
            Wvref.en=1'b1;
            Wvref.value=0.0;
`else
            vref = 0;
`endif    
      end
   end 
   else begin
`ifdef WPIN_UART_EN
         Wvref.en=1'b0;
`else 
      vref= 1'bx;
`endif
   end
end


endmodule
`endif //SYNTHESIS
