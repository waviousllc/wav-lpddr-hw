/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
*****************************************************************************
*
* Module    : ddr_dq_drvr_lpbk_wrapper.sv
* Date      : 2020-04-19
* Desciption: DQ Driver with loopback
* Author    : shadzibabic
*
****************************************************************************/

`include "ddr_global_define.vh"
`include "ddr_project_define.vh"
`include "ddr_dq_drvr_lpbk_wrapper_define.vh"
`include "ddr_dq_drvr_lpbk_wrapper_cmn_define.vh"

import ddr_global_pkg::*;

module ddr_dq_drvr_lpbk_wrapper #(
   parameter P0WIDTH = 6,
   parameter P1WIDTH = 19
)
(
   input  logic [P0WIDTH-1:0] i_drvr_cfg,
   input  logic [P1WIDTH-1:0] i_drvr_cmn_cfg,
   input  logic i_freeze_n,
   input  logic i_hiz_n,
   input  logic i_d_n,
   input  logic i_oe,
   input  logic i_bs_mode_n,
   input  logic i_bs_oe,
   input  logic i_bs_ie,
   input  logic i_d_bs,
   inout  wire  pad,
   output wire  o_d_lpbk,
   output wire  o_rx_in
);

`ifndef WLOGIC_NO_PG
   wire vdda, vdd_aon, vddq, vss;
   assign vdda    = 1'b1;
   assign vdd_aon = 1'b1;
   assign vddq    = 1'b1;
   assign vss     = 1'b0;
`endif

   logic lpbk_ena;
`ifndef DDR_IO_WRAPPER_BEHAV
   ddr_wcm_mux #(.DWIDTH(1)) u_mux_lpbk_ena (.i_sel(i_bs_mode_n), .i_a(i_bs_ie), .i_b(i_drvr_cmn_cfg[`DDR_ANA_DQ_DRVR_LPBK_LPBK_EN_FIELD]), .o_z(lpbk_ena));
`else
   assign lpbk_ena =  i_bs_mode_n ? i_drvr_cmn_cfg[`DDR_ANA_DQ_DRVR_LPBK_LPBK_EN_FIELD] : i_bs_ie;
`endif

   logic bs_ena;
`ifndef DDR_IO_WRAPPER_BEHAV
   ddr_wcm_mux #(.DWIDTH(1)) u_mux_bs_ena (.i_sel(i_bs_mode_n), .i_a(i_bs_oe), .i_b(i_drvr_cmn_cfg[`DDR_ANA_DQ_DRVR_LPBK_BS_EN_FIELD]), .o_z(bs_ena));
`else
   assign bs_ena   =  i_bs_mode_n ? i_drvr_cmn_cfg[`DDR_ANA_DQ_DRVR_LPBK_BS_EN_FIELD]   : i_bs_oe;
`endif

   // See wphy_lp4x5_dq_drv.doc, section 1.7.1 for details on driver configuration
   // for freeze and hiz ...
   //   if (freeze)   {d_drv_impd, d_ovrd, d_ovrd_val} = {2’h1, 3’h1, 1’b0}
   //   else if (hiz) {d_drv_impd, d_ovrd, d_ovrd_val} = {2’h0, 3’h1, 1’b0}

   logic [2:0] ovrd;
   // See wphy_lp4x5_dq_drv.doc, section 1.7.1 for details on driver configuration
`ifndef DDR_IO_WRAPPER_BEHAV
   logic [2:0] lpbk_ovrd_sel_oe;
   logic [2:0] oe_bus_b;
   logic [2:0] ovrd_mux_1;
   logic [2:0] ovrd_mux_2;
   logic [2:0] ovrd_mux_3;

   ddr_wcm_inv u_inv_oe_int_0  ( .i_a(i_oe), .o_z(oe_bus_b[0]));
   ddr_wcm_inv u_inv_oe_int_1  ( .i_a(i_oe), .o_z(oe_bus_b[1]));
   ddr_wcm_inv u_inv_oe_int_2  ( .i_a(i_oe), .o_z(oe_bus_b[2]));

  //TODO - add tiehi/lo
   ddr_wcm_and #(3) u_and_ovrd_oe ( .i_a(oe_bus_b), .i_b(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_OVRD_SEL_FIELD]), .o_z(lpbk_ovrd_sel_oe));
   ddr_wcm_mux #(3) u_mux_ovrd_1 (.i_sel(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_SW_OVR_FIELD]), .i_a(lpbk_ovrd_sel_oe), .i_b(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_OVRD_SEL_FIELD]), .o_z(ovrd_mux_1));
   ddr_wcm_mux #(3) u_mux_ovrd_2 (.i_sel(i_bs_mode_n), .i_a(3'h1), .i_b(ovrd_mux_1), .o_z(ovrd_mux_2));
   ddr_wcm_mux #(3) u_mux_ovrd_3 (.i_sel(i_hiz_n), .i_a(3'h1), .i_b(ovrd_mux_2), .o_z(ovrd_mux_3));
   ddr_wcm_mux #(3) u_mux_ovrd_4 (.i_sel(i_freeze_n), .i_a(3'h1), .i_b(ovrd_mux_3), .o_z(ovrd));
`else
   assign ovrd = i_freeze_n ? i_hiz_n ? i_bs_mode_n ?
                    i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_SW_OVR_FIELD] ?
                    i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_OVRD_SEL_FIELD] :
                    {3{~i_oe}} & i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_OVRD_SEL_FIELD]
                 : 3'h1 : 3'h1 : 3'h1;
`endif

   logic [2:0] impd;
`ifndef DDR_IO_WRAPPER_BEHAV
   logic lpbk_sw_ovrd;
   logic [2:0] oe_bus;
   logic [2:0] impd_mux_1;
   logic [2:0] impd_mux_2;
   logic [2:0] impd_mux_3;

   //assign oe_bus[0] = oe;
   //assign oe_bus[1] = oe;
   //assign oe_bus[2] = oe;

  //TODO - add tiehi/lo
   ddr_wcm_or   u_or_sw_ovrd (.i_a(i_oe), .i_b(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_SW_OVR_FIELD]), .o_z(lpbk_sw_ovrd));
   ddr_wcm_mux #(.DWIDTH(3)) u_mux_impd_1 (.i_sel(lpbk_sw_ovrd), .i_a(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_RX_IMPD_FIELD]), .i_b(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_TX_IMPD_FIELD]), .o_z(impd_mux_1));
   ddr_wcm_mux #(.DWIDTH(3)) u_mux_impd_2 (.i_sel(i_bs_mode_n), .i_a(3'h0), .i_b(impd_mux_1), .o_z(impd_mux_2));
   ddr_wcm_mux #(.DWIDTH(3)) u_mux_impd_3 (.i_sel(i_hiz_n), .i_a(3'h0), .i_b(impd_mux_2), .o_z(impd_mux_3));
   ddr_wcm_mux #(.DWIDTH(3)) u_mux_impd_4 (.i_sel(i_freeze_n), .i_a(3'h1), .i_b(impd_mux_3), .o_z(impd));
`else
   assign impd = i_freeze_n ? i_hiz_n ? i_bs_mode_n ?
                    i_oe | i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_SW_OVR_FIELD] ?
                    i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_TX_IMPD_FIELD]:
                    i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_RX_IMPD_FIELD]
                 : 3'h0 : 3'h0 : 3'h1;
`endif

   logic ovrd_val;
`ifndef DDR_IO_WRAPPER_BEHAV
   logic  val_mux_1;
   logic  val_mux_2;
   logic  val_mux_3;

  //TODO - add tiehi/lo
   ddr_wcm_mux  u_mux_val_1 (.i_sel(i_bs_mode_n), .i_a(1'h0), .i_b(i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_OVRD_VAL_FIELD]), .o_z(val_mux_1));
   ddr_wcm_mux  u_mux_val_2 (.i_sel(i_hiz_n), .i_a(1'h0), .i_b(val_mux_1), .o_z(val_mux_2));
   ddr_wcm_mux  u_mux_val_3 (.i_sel(i_freeze_n), .i_a(1'h0), .i_b(val_mux_2), .o_z(ovrd_val));
`else
   assign ovrd_val = i_freeze_n ? i_hiz_n ? i_bs_mode_n ?
                    i_drvr_cfg[`DDR_ANA_DQ_DRVR_LPBK_OVRD_VAL_FIELD]
                 : 1'h0 : 1'h0 : 1'h0;
`endif

   wphy_lp4x5_dq_drvr_w_lpbk u_dq_drvr_w_lpbk (
      .pad           (pad),
      //.d_in          (i_d),
      .d_in_c          (i_d_n),
      .d_bs_din      (i_d_bs),
      .d_bs_ena      (bs_ena),
      .d_lpbk_ena    (lpbk_ena),
      .freeze_n      (i_freeze_n),
      .d_lpbk_out    (o_d_lpbk),
      .rx_in         (o_rx_in),
      .d_ovrd        (ovrd),
      .d_ovrd_val    (ovrd_val),
      .d_drv_impd    (impd),
      .d_ncal        (i_drvr_cmn_cfg[`DDR_ANA_DQ_DRVR_LPBK_NCAL_FIELD]),
      .d_pcal        (i_drvr_cmn_cfg[`DDR_ANA_DQ_DRVR_LPBK_PCAL_FIELD])
`ifndef WLOGIC_NO_PG
      ,.vdda         (vdda),
      .vdd_aon       (vdd_aon),
      .vddq          (vddq),
      .vss           (vss)
`endif
   );

endmodule
