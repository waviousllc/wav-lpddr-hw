
/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`include "ddr_global_define.vh"
`include "ddr_project_define.vh"
`include "ddr_dq_csr_defs.vh"

import ddr_global_pkg::*;

module ddr_dq_ahb_csr #(
   parameter AWIDTH = 32,
   parameter DWIDTH = 32
) (

   input   logic                i_hclk,
   input   logic                i_hreset,
   input   logic [AWIDTH-1:0]   i_haddr,
   input   logic                i_hwrite,
   input   logic                i_hsel,
   input   logic [DWIDTH-1:0]   i_hwdata,
   input   logic [1:0]          i_htrans,
   input   logic [2:0]          i_hsize,
   input   logic [2:0]          i_hburst,
   input   logic                i_hreadyin,
   output  logic                o_hready,
   output  logic [DWIDTH-1:0]   o_hrdata,
   output  logic [1:0]          o_hresp,
   output  logic [`DDR_DQ_TOP_CFG_RANGE] o_dq_top_cfg,
   input   logic [`DDR_DQ_TOP_STA_RANGE] i_dq_top_sta,
   input   logic [`DDR_DQ_DQ_RX_BSCAN_STA_RANGE] i_dq_dq_rx_bscan_sta,
   output  logic [`DDR_DQ_DQ_RX_M0_CFG_RANGE] o_dq_dq_rx_m0_cfg,
   output  logic [`DDR_DQ_DQ_RX_M1_CFG_RANGE] o_dq_dq_rx_m1_cfg,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_0_RANGE] o_dq_dq_rx_io_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_1_RANGE] o_dq_dq_rx_io_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_2_RANGE] o_dq_dq_rx_io_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_3_RANGE] o_dq_dq_rx_io_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_4_RANGE] o_dq_dq_rx_io_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_5_RANGE] o_dq_dq_rx_io_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_6_RANGE] o_dq_dq_rx_io_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_7_RANGE] o_dq_dq_rx_io_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R0_CFG_8_RANGE] o_dq_dq_rx_io_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_0_RANGE] o_dq_dq_rx_io_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_1_RANGE] o_dq_dq_rx_io_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_2_RANGE] o_dq_dq_rx_io_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_3_RANGE] o_dq_dq_rx_io_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_4_RANGE] o_dq_dq_rx_io_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_5_RANGE] o_dq_dq_rx_io_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_6_RANGE] o_dq_dq_rx_io_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_7_RANGE] o_dq_dq_rx_io_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_IO_M0_R1_CFG_8_RANGE] o_dq_dq_rx_io_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_0_RANGE] o_dq_dq_rx_io_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_1_RANGE] o_dq_dq_rx_io_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_2_RANGE] o_dq_dq_rx_io_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_3_RANGE] o_dq_dq_rx_io_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_4_RANGE] o_dq_dq_rx_io_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_5_RANGE] o_dq_dq_rx_io_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_6_RANGE] o_dq_dq_rx_io_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_7_RANGE] o_dq_dq_rx_io_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R0_CFG_8_RANGE] o_dq_dq_rx_io_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_0_RANGE] o_dq_dq_rx_io_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_1_RANGE] o_dq_dq_rx_io_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_2_RANGE] o_dq_dq_rx_io_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_3_RANGE] o_dq_dq_rx_io_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_4_RANGE] o_dq_dq_rx_io_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_5_RANGE] o_dq_dq_rx_io_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_6_RANGE] o_dq_dq_rx_io_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_7_RANGE] o_dq_dq_rx_io_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_IO_M1_R1_CFG_8_RANGE] o_dq_dq_rx_io_m1_r1_cfg_8,
   input   logic [`DDR_DQ_DQ_RX_IO_STA_RANGE] i_dq_dq_rx_io_sta,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_0_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_1_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_2_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_3_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_4_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_5_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_6_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_7_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R0_CFG_8_RANGE] o_dq_dq_rx_sa_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_0_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_1_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_2_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_3_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_4_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_5_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_6_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_7_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_M0_R1_CFG_8_RANGE] o_dq_dq_rx_sa_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_0_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_1_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_2_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_3_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_4_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_5_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_6_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_7_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R0_CFG_8_RANGE] o_dq_dq_rx_sa_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_0_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_1_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_2_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_3_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_4_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_5_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_6_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_7_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_M1_R1_CFG_8_RANGE] o_dq_dq_rx_sa_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_0_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_1_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_2_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_3_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_4_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_5_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_6_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_7_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R0_CFG_8_RANGE] o_dq_dq_rx_sa_dly_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_0_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_1_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_2_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_3_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_4_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_5_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_6_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_7_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M0_R1_CFG_8_RANGE] o_dq_dq_rx_sa_dly_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_0_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_1_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_2_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_3_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_4_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_5_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_6_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_7_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R0_CFG_8_RANGE] o_dq_dq_rx_sa_dly_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_0_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_1_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_2_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_3_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_4_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_5_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_6_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_7_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_RX_SA_DLY_M1_R1_CFG_8_RANGE] o_dq_dq_rx_sa_dly_m1_r1_cfg_8,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_0_RANGE] i_dq_dq_rx_sa_sta_0,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_1_RANGE] i_dq_dq_rx_sa_sta_1,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_2_RANGE] i_dq_dq_rx_sa_sta_2,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_3_RANGE] i_dq_dq_rx_sa_sta_3,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_4_RANGE] i_dq_dq_rx_sa_sta_4,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_5_RANGE] i_dq_dq_rx_sa_sta_5,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_6_RANGE] i_dq_dq_rx_sa_sta_6,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_7_RANGE] i_dq_dq_rx_sa_sta_7,
   input   logic [`DDR_DQ_DQ_RX_SA_STA_8_RANGE] i_dq_dq_rx_sa_sta_8,
   output  logic [`DDR_DQ_DQ_TX_BSCAN_CFG_RANGE] o_dq_dq_tx_bscan_cfg,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_0_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_1_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_2_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_3_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_4_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_5_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_6_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_7_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M0_CFG_8_RANGE] o_dq_dq_tx_egress_ana_m0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_0_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_1_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_2_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_3_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_4_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_5_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_6_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_7_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_ANA_M1_CFG_8_RANGE] o_dq_dq_tx_egress_ana_m1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_0_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_1_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_2_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_3_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_4_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_5_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_6_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_7_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M0_CFG_8_RANGE] o_dq_dq_tx_egress_dig_m0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_0_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_1_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_2_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_3_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_4_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_5_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_6_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_7_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_EGRESS_DIG_M1_CFG_8_RANGE] o_dq_dq_tx_egress_dig_m1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_ODR_PI_M0_R0_CFG_RANGE] o_dq_dq_tx_odr_pi_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_ODR_PI_M0_R1_CFG_RANGE] o_dq_dq_tx_odr_pi_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_ODR_PI_M1_R0_CFG_RANGE] o_dq_dq_tx_odr_pi_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_ODR_PI_M1_R1_CFG_RANGE] o_dq_dq_tx_odr_pi_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_0_M0_R0_CFG_RANGE] o_dq_dq_tx_qdr_pi_0_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_0_M0_R1_CFG_RANGE] o_dq_dq_tx_qdr_pi_0_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_0_M1_R0_CFG_RANGE] o_dq_dq_tx_qdr_pi_0_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_0_M1_R1_CFG_RANGE] o_dq_dq_tx_qdr_pi_0_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_1_M0_R0_CFG_RANGE] o_dq_dq_tx_qdr_pi_1_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_1_M0_R1_CFG_RANGE] o_dq_dq_tx_qdr_pi_1_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_1_M1_R0_CFG_RANGE] o_dq_dq_tx_qdr_pi_1_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_QDR_PI_1_M1_R1_CFG_RANGE] o_dq_dq_tx_qdr_pi_1_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_0_M0_R0_CFG_RANGE] o_dq_dq_tx_ddr_pi_0_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_0_M0_R1_CFG_RANGE] o_dq_dq_tx_ddr_pi_0_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_0_M1_R0_CFG_RANGE] o_dq_dq_tx_ddr_pi_0_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_0_M1_R1_CFG_RANGE] o_dq_dq_tx_ddr_pi_0_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_1_M0_R0_CFG_RANGE] o_dq_dq_tx_ddr_pi_1_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_1_M0_R1_CFG_RANGE] o_dq_dq_tx_ddr_pi_1_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_1_M1_R0_CFG_RANGE] o_dq_dq_tx_ddr_pi_1_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_DDR_PI_1_M1_R1_CFG_RANGE] o_dq_dq_tx_ddr_pi_1_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_PI_RT_M0_R0_CFG_RANGE] o_dq_dq_tx_pi_rt_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_PI_RT_M0_R1_CFG_RANGE] o_dq_dq_tx_pi_rt_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_PI_RT_M1_R0_CFG_RANGE] o_dq_dq_tx_pi_rt_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_PI_RT_M1_R1_CFG_RANGE] o_dq_dq_tx_pi_rt_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_RT_M0_R0_CFG_RANGE] o_dq_dq_tx_rt_m0_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_RT_M0_R1_CFG_RANGE] o_dq_dq_tx_rt_m0_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_RT_M1_R0_CFG_RANGE] o_dq_dq_tx_rt_m1_r0_cfg,
   output  logic [`DDR_DQ_DQ_TX_RT_M1_R1_CFG_RANGE] o_dq_dq_tx_rt_m1_r1_cfg,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_0_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_1_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_2_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_3_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_4_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_5_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_6_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_7_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R0_CFG_8_RANGE] o_dq_dq_tx_sdr_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_0_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_1_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_2_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_3_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_4_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_5_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_6_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_7_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_M0_R1_CFG_8_RANGE] o_dq_dq_tx_sdr_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_0_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_1_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_2_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_3_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_4_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_5_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_6_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_7_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R0_CFG_8_RANGE] o_dq_dq_tx_sdr_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_0_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_1_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_2_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_3_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_4_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_5_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_6_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_7_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_M1_R1_CFG_8_RANGE] o_dq_dq_tx_sdr_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_RANGE] o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_RANGE] o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_RANGE] o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_RANGE] o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_0_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_1_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_2_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_3_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_4_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_5_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_6_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_7_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R0_CFG_8_RANGE] o_dq_dq_tx_ddr_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_0_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_1_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_2_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_3_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_4_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_5_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_6_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_7_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_M0_R1_CFG_8_RANGE] o_dq_dq_tx_ddr_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_0_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_1_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_2_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_3_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_4_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_5_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_6_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_7_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R0_CFG_8_RANGE] o_dq_dq_tx_ddr_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_0_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_1_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_2_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_3_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_4_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_5_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_6_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_7_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_M1_R1_CFG_8_RANGE] o_dq_dq_tx_ddr_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_RANGE] o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_RANGE] o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_0_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_1_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_2_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_3_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_4_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_5_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_6_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_7_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R0_CFG_8_RANGE] o_dq_dq_tx_qdr_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_0_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_1_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_2_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_3_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_4_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_5_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_6_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_7_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_M0_R1_CFG_8_RANGE] o_dq_dq_tx_qdr_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_0_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_1_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_2_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_3_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_4_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_5_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_6_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_7_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R0_CFG_8_RANGE] o_dq_dq_tx_qdr_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_0_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_1_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_2_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_3_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_4_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_5_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_6_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_7_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_M1_R1_CFG_8_RANGE] o_dq_dq_tx_qdr_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_RANGE] o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_RANGE] o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_0_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_1_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_2_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_3_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_4_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_5_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_6_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_7_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R0_CFG_8_RANGE] o_dq_dq_tx_lpde_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_0_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_1_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_2_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_3_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_4_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_5_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_6_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_7_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M0_R1_CFG_8_RANGE] o_dq_dq_tx_lpde_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_0_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_1_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_2_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_3_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_4_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_5_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_6_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_7_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R0_CFG_8_RANGE] o_dq_dq_tx_lpde_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_0_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_1_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_2_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_3_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_4_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_5_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_6_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_7_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_LPDE_M1_R1_CFG_8_RANGE] o_dq_dq_tx_lpde_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_0_RANGE] o_dq_dq_tx_io_m0_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_1_RANGE] o_dq_dq_tx_io_m0_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_2_RANGE] o_dq_dq_tx_io_m0_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_3_RANGE] o_dq_dq_tx_io_m0_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_4_RANGE] o_dq_dq_tx_io_m0_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_5_RANGE] o_dq_dq_tx_io_m0_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_6_RANGE] o_dq_dq_tx_io_m0_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_7_RANGE] o_dq_dq_tx_io_m0_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_IO_M0_CFG_8_RANGE] o_dq_dq_tx_io_m0_cfg_8,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_0_RANGE] o_dq_dq_tx_io_m1_cfg_0,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_1_RANGE] o_dq_dq_tx_io_m1_cfg_1,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_2_RANGE] o_dq_dq_tx_io_m1_cfg_2,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_3_RANGE] o_dq_dq_tx_io_m1_cfg_3,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_4_RANGE] o_dq_dq_tx_io_m1_cfg_4,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_5_RANGE] o_dq_dq_tx_io_m1_cfg_5,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_6_RANGE] o_dq_dq_tx_io_m1_cfg_6,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_7_RANGE] o_dq_dq_tx_io_m1_cfg_7,
   output  logic [`DDR_DQ_DQ_TX_IO_M1_CFG_8_RANGE] o_dq_dq_tx_io_m1_cfg_8,
   output  logic [`DDR_DQ_DQS_RX_M0_CFG_RANGE] o_dq_dqs_rx_m0_cfg,
   output  logic [`DDR_DQ_DQS_RX_M1_CFG_RANGE] o_dq_dqs_rx_m1_cfg,
   input   logic [`DDR_DQ_DQS_RX_BSCAN_STA_RANGE] i_dq_dqs_rx_bscan_sta,
   output  logic [`DDR_DQ_DQS_RX_SDR_LPDE_M0_R0_CFG_RANGE] o_dq_dqs_rx_sdr_lpde_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_SDR_LPDE_M0_R1_CFG_RANGE] o_dq_dqs_rx_sdr_lpde_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_SDR_LPDE_M1_R0_CFG_RANGE] o_dq_dqs_rx_sdr_lpde_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_SDR_LPDE_M1_R1_CFG_RANGE] o_dq_dqs_rx_sdr_lpde_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_REN_PI_M0_R0_CFG_RANGE] o_dq_dqs_rx_ren_pi_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_REN_PI_M0_R1_CFG_RANGE] o_dq_dqs_rx_ren_pi_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_REN_PI_M1_R0_CFG_RANGE] o_dq_dqs_rx_ren_pi_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_REN_PI_M1_R1_CFG_RANGE] o_dq_dqs_rx_ren_pi_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_RCS_PI_M0_R0_CFG_RANGE] o_dq_dqs_rx_rcs_pi_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_RCS_PI_M0_R1_CFG_RANGE] o_dq_dqs_rx_rcs_pi_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_RCS_PI_M1_R0_CFG_RANGE] o_dq_dqs_rx_rcs_pi_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_RCS_PI_M1_R1_CFG_RANGE] o_dq_dqs_rx_rcs_pi_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_0_M0_R0_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_0_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_0_M0_R1_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_0_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_0_M1_R0_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_0_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_0_M1_R1_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_0_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_1_M0_R0_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_1_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_1_M0_R1_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_1_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_1_M1_R0_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_1_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_RDQS_PI_1_M1_R1_CFG_RANGE] o_dq_dqs_rx_rdqs_pi_1_m1_r1_cfg,
   input   logic [`DDR_DQ_DQS_RX_PI_STA_RANGE] i_dq_dqs_rx_pi_sta,
   output  logic [`DDR_DQ_DQS_RX_IO_M0_R0_CFG_0_RANGE] o_dq_dqs_rx_io_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_IO_M0_R0_CFG_1_RANGE] o_dq_dqs_rx_io_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_IO_M0_R1_CFG_0_RANGE] o_dq_dqs_rx_io_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_IO_M0_R1_CFG_1_RANGE] o_dq_dqs_rx_io_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_IO_M1_R0_CFG_0_RANGE] o_dq_dqs_rx_io_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_IO_M1_R0_CFG_1_RANGE] o_dq_dqs_rx_io_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_IO_M1_R1_CFG_0_RANGE] o_dq_dqs_rx_io_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_IO_M1_R1_CFG_1_RANGE] o_dq_dqs_rx_io_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_IO_CMN_M0_R0_CFG_RANGE] o_dq_dqs_rx_io_cmn_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_IO_CMN_M0_R1_CFG_RANGE] o_dq_dqs_rx_io_cmn_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_RX_IO_CMN_M1_R0_CFG_RANGE] o_dq_dqs_rx_io_cmn_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_RX_IO_CMN_M1_R1_CFG_RANGE] o_dq_dqs_rx_io_cmn_m1_r1_cfg,
   input   logic [`DDR_DQ_DQS_RX_IO_STA_RANGE] i_dq_dqs_rx_io_sta,
   output  logic [`DDR_DQ_DQS_RX_SA_M0_R0_CFG_0_RANGE] o_dq_dqs_rx_sa_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_SA_M0_R0_CFG_1_RANGE] o_dq_dqs_rx_sa_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_SA_M0_R1_CFG_0_RANGE] o_dq_dqs_rx_sa_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_SA_M0_R1_CFG_1_RANGE] o_dq_dqs_rx_sa_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_SA_M1_R0_CFG_0_RANGE] o_dq_dqs_rx_sa_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_SA_M1_R0_CFG_1_RANGE] o_dq_dqs_rx_sa_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_SA_M1_R1_CFG_0_RANGE] o_dq_dqs_rx_sa_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_RX_SA_M1_R1_CFG_1_RANGE] o_dq_dqs_rx_sa_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_RX_SA_CMN_CFG_RANGE] o_dq_dqs_rx_sa_cmn_cfg,
   output  logic [`DDR_DQ_DQS_TX_M0_CFG_RANGE] o_dq_dqs_tx_m0_cfg,
   output  logic [`DDR_DQ_DQS_TX_M1_CFG_RANGE] o_dq_dqs_tx_m1_cfg,
   output  logic [`DDR_DQ_DQS_TX_BSCAN_CTRL_CFG_RANGE] o_dq_dqs_tx_bscan_ctrl_cfg,
   output  logic [`DDR_DQ_DQS_TX_BSCAN_CFG_RANGE] o_dq_dqs_tx_bscan_cfg,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_0_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_1_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_2_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_3_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_4_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_5_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_6_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_7_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M0_CFG_8_RANGE] o_dq_dqs_tx_egress_ana_m0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_0_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_1_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_2_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_3_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_4_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_5_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_6_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_7_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_ANA_M1_CFG_8_RANGE] o_dq_dqs_tx_egress_ana_m1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_0_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_1_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_2_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_3_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_4_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_5_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_6_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_7_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M0_CFG_8_RANGE] o_dq_dqs_tx_egress_dig_m0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_0_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_1_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_2_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_3_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_4_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_5_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_6_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_7_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_EGRESS_DIG_M1_CFG_8_RANGE] o_dq_dqs_tx_egress_dig_m1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_ODR_PI_M0_R0_CFG_RANGE] o_dq_dqs_tx_odr_pi_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_ODR_PI_M0_R1_CFG_RANGE] o_dq_dqs_tx_odr_pi_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_ODR_PI_M1_R0_CFG_RANGE] o_dq_dqs_tx_odr_pi_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_ODR_PI_M1_R1_CFG_RANGE] o_dq_dqs_tx_odr_pi_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_0_M0_R0_CFG_RANGE] o_dq_dqs_tx_qdr_pi_0_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_0_M0_R1_CFG_RANGE] o_dq_dqs_tx_qdr_pi_0_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_0_M1_R0_CFG_RANGE] o_dq_dqs_tx_qdr_pi_0_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_0_M1_R1_CFG_RANGE] o_dq_dqs_tx_qdr_pi_0_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_1_M0_R0_CFG_RANGE] o_dq_dqs_tx_qdr_pi_1_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_1_M0_R1_CFG_RANGE] o_dq_dqs_tx_qdr_pi_1_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_1_M1_R0_CFG_RANGE] o_dq_dqs_tx_qdr_pi_1_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_QDR_PI_1_M1_R1_CFG_RANGE] o_dq_dqs_tx_qdr_pi_1_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_0_M0_R0_CFG_RANGE] o_dq_dqs_tx_ddr_pi_0_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_0_M0_R1_CFG_RANGE] o_dq_dqs_tx_ddr_pi_0_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_0_M1_R0_CFG_RANGE] o_dq_dqs_tx_ddr_pi_0_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_0_M1_R1_CFG_RANGE] o_dq_dqs_tx_ddr_pi_0_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_1_M0_R0_CFG_RANGE] o_dq_dqs_tx_ddr_pi_1_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_1_M0_R1_CFG_RANGE] o_dq_dqs_tx_ddr_pi_1_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_1_M1_R0_CFG_RANGE] o_dq_dqs_tx_ddr_pi_1_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_DDR_PI_1_M1_R1_CFG_RANGE] o_dq_dqs_tx_ddr_pi_1_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_PI_RT_M0_R0_CFG_RANGE] o_dq_dqs_tx_pi_rt_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_PI_RT_M0_R1_CFG_RANGE] o_dq_dqs_tx_pi_rt_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_PI_RT_M1_R0_CFG_RANGE] o_dq_dqs_tx_pi_rt_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_PI_RT_M1_R1_CFG_RANGE] o_dq_dqs_tx_pi_rt_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_SDR_PI_M0_R0_CFG_RANGE] o_dq_dqs_tx_sdr_pi_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_SDR_PI_M0_R1_CFG_RANGE] o_dq_dqs_tx_sdr_pi_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_SDR_PI_M1_R0_CFG_RANGE] o_dq_dqs_tx_sdr_pi_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_SDR_PI_M1_R1_CFG_RANGE] o_dq_dqs_tx_sdr_pi_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_DFI_PI_M0_R0_CFG_RANGE] o_dq_dqs_tx_dfi_pi_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_DFI_PI_M0_R1_CFG_RANGE] o_dq_dqs_tx_dfi_pi_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_DFI_PI_M1_R0_CFG_RANGE] o_dq_dqs_tx_dfi_pi_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_DFI_PI_M1_R1_CFG_RANGE] o_dq_dqs_tx_dfi_pi_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_RT_M0_R0_CFG_RANGE] o_dq_dqs_tx_rt_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_RT_M0_R1_CFG_RANGE] o_dq_dqs_tx_rt_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_RT_M1_R0_CFG_RANGE] o_dq_dqs_tx_rt_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_RT_M1_R1_CFG_RANGE] o_dq_dqs_tx_rt_m1_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_sdr_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_sdr_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_sdr_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_sdr_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_X_SEL_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_ddr_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_ddr_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_ddr_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_ddr_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_DDR_X_SEL_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_qdr_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_qdr_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_qdr_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_qdr_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_2_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_3_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_4_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_5_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_6_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_7_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R0_CFG_8_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_2_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_3_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_4_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_5_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_6_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_7_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M0_R1_CFG_8_RANGE] o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_2_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_3_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_4_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_5_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_6_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_7_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R0_CFG_8_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_2_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_2,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_3_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_3,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_4_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_4,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_5_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_5,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_6_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_6,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_7_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_7,
   output  logic [`DDR_DQ_DQS_TX_QDR_X_SEL_M1_R1_CFG_8_RANGE] o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_8,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M0_R0_CFG_0_RANGE] o_dq_dqs_tx_lpde_m0_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M0_R0_CFG_1_RANGE] o_dq_dqs_tx_lpde_m0_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M0_R1_CFG_0_RANGE] o_dq_dqs_tx_lpde_m0_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M0_R1_CFG_1_RANGE] o_dq_dqs_tx_lpde_m0_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M1_R0_CFG_0_RANGE] o_dq_dqs_tx_lpde_m1_r0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M1_R0_CFG_1_RANGE] o_dq_dqs_tx_lpde_m1_r0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M1_R1_CFG_0_RANGE] o_dq_dqs_tx_lpde_m1_r1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_LPDE_M1_R1_CFG_1_RANGE] o_dq_dqs_tx_lpde_m1_r1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_IO_M0_CFG_0_RANGE] o_dq_dqs_tx_io_m0_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_IO_M0_CFG_1_RANGE] o_dq_dqs_tx_io_m0_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_IO_M1_CFG_0_RANGE] o_dq_dqs_tx_io_m1_cfg_0,
   output  logic [`DDR_DQ_DQS_TX_IO_M1_CFG_1_RANGE] o_dq_dqs_tx_io_m1_cfg_1,
   output  logic [`DDR_DQ_DQS_TX_IO_CMN_M0_R0_CFG_RANGE] o_dq_dqs_tx_io_cmn_m0_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_IO_CMN_M0_R1_CFG_RANGE] o_dq_dqs_tx_io_cmn_m0_r1_cfg,
   output  logic [`DDR_DQ_DQS_TX_IO_CMN_M1_R0_CFG_RANGE] o_dq_dqs_tx_io_cmn_m1_r0_cfg,
   output  logic [`DDR_DQ_DQS_TX_IO_CMN_M1_R1_CFG_RANGE] o_dq_dqs_tx_io_cmn_m1_r1_cfg
);

   logic                slv_write;
   logic                slv_read;
   logic                slv_error;
   logic [AWIDTH-1:0]   slv_addr;
   logic [DWIDTH-1:0]   slv_wdata;
   logic [DWIDTH-1:0]   slv_rdata;
   logic                slv_ready;

   ddr_ahb_slave #(
      .AWIDTH(AWIDTH),
      .DWIDTH(DWIDTH)
   ) ahb_slave (
      .i_hclk     (i_hclk),
      .i_hreset   (i_hreset),
      .i_haddr    (i_haddr),
      .i_hwrite   (i_hwrite),
      .i_hsel     (i_hsel),
      .i_hwdata   (i_hwdata),
      .i_htrans   (i_htrans),
      .i_hsize    (i_hsize),
      .i_hburst   (i_hburst),
      .i_hreadyin (i_hreadyin),
      .o_hready   (o_hready),
      .o_hrdata   (o_hrdata),
      .o_hresp    (o_hresp),
      .o_write    (slv_write),
      .o_read     (slv_read),
      .o_wdata    (slv_wdata),
      .o_addr     (slv_addr),
      .i_rdata    (slv_rdata),
      .i_error    (slv_error),
      .i_ready    (slv_ready)
   );

   ddr_dq_csr #(
      .AWIDTH(AWIDTH),
      .DWIDTH(DWIDTH)
   ) dq_csr (
      .i_hclk   (i_hclk),
      .i_hreset (i_hreset),
      .i_write  (slv_write),
      .i_read   (slv_read),
      .i_wdata  (slv_wdata),
      .i_addr   (slv_addr),
      .o_rdata  (slv_rdata),
      .o_error  (slv_error),
      .o_ready  (slv_ready),
      .o_dq_top_cfg (o_dq_top_cfg),
      .i_dq_top_sta (i_dq_top_sta),
      .i_dq_dq_rx_bscan_sta (i_dq_dq_rx_bscan_sta),
      .o_dq_dq_rx_m0_cfg (o_dq_dq_rx_m0_cfg),
      .o_dq_dq_rx_m1_cfg (o_dq_dq_rx_m1_cfg),
      .o_dq_dq_rx_io_m0_r0_cfg_0 (o_dq_dq_rx_io_m0_r0_cfg_0),
      .o_dq_dq_rx_io_m0_r0_cfg_1 (o_dq_dq_rx_io_m0_r0_cfg_1),
      .o_dq_dq_rx_io_m0_r0_cfg_2 (o_dq_dq_rx_io_m0_r0_cfg_2),
      .o_dq_dq_rx_io_m0_r0_cfg_3 (o_dq_dq_rx_io_m0_r0_cfg_3),
      .o_dq_dq_rx_io_m0_r0_cfg_4 (o_dq_dq_rx_io_m0_r0_cfg_4),
      .o_dq_dq_rx_io_m0_r0_cfg_5 (o_dq_dq_rx_io_m0_r0_cfg_5),
      .o_dq_dq_rx_io_m0_r0_cfg_6 (o_dq_dq_rx_io_m0_r0_cfg_6),
      .o_dq_dq_rx_io_m0_r0_cfg_7 (o_dq_dq_rx_io_m0_r0_cfg_7),
      .o_dq_dq_rx_io_m0_r0_cfg_8 (o_dq_dq_rx_io_m0_r0_cfg_8),
      .o_dq_dq_rx_io_m0_r1_cfg_0 (o_dq_dq_rx_io_m0_r1_cfg_0),
      .o_dq_dq_rx_io_m0_r1_cfg_1 (o_dq_dq_rx_io_m0_r1_cfg_1),
      .o_dq_dq_rx_io_m0_r1_cfg_2 (o_dq_dq_rx_io_m0_r1_cfg_2),
      .o_dq_dq_rx_io_m0_r1_cfg_3 (o_dq_dq_rx_io_m0_r1_cfg_3),
      .o_dq_dq_rx_io_m0_r1_cfg_4 (o_dq_dq_rx_io_m0_r1_cfg_4),
      .o_dq_dq_rx_io_m0_r1_cfg_5 (o_dq_dq_rx_io_m0_r1_cfg_5),
      .o_dq_dq_rx_io_m0_r1_cfg_6 (o_dq_dq_rx_io_m0_r1_cfg_6),
      .o_dq_dq_rx_io_m0_r1_cfg_7 (o_dq_dq_rx_io_m0_r1_cfg_7),
      .o_dq_dq_rx_io_m0_r1_cfg_8 (o_dq_dq_rx_io_m0_r1_cfg_8),
      .o_dq_dq_rx_io_m1_r0_cfg_0 (o_dq_dq_rx_io_m1_r0_cfg_0),
      .o_dq_dq_rx_io_m1_r0_cfg_1 (o_dq_dq_rx_io_m1_r0_cfg_1),
      .o_dq_dq_rx_io_m1_r0_cfg_2 (o_dq_dq_rx_io_m1_r0_cfg_2),
      .o_dq_dq_rx_io_m1_r0_cfg_3 (o_dq_dq_rx_io_m1_r0_cfg_3),
      .o_dq_dq_rx_io_m1_r0_cfg_4 (o_dq_dq_rx_io_m1_r0_cfg_4),
      .o_dq_dq_rx_io_m1_r0_cfg_5 (o_dq_dq_rx_io_m1_r0_cfg_5),
      .o_dq_dq_rx_io_m1_r0_cfg_6 (o_dq_dq_rx_io_m1_r0_cfg_6),
      .o_dq_dq_rx_io_m1_r0_cfg_7 (o_dq_dq_rx_io_m1_r0_cfg_7),
      .o_dq_dq_rx_io_m1_r0_cfg_8 (o_dq_dq_rx_io_m1_r0_cfg_8),
      .o_dq_dq_rx_io_m1_r1_cfg_0 (o_dq_dq_rx_io_m1_r1_cfg_0),
      .o_dq_dq_rx_io_m1_r1_cfg_1 (o_dq_dq_rx_io_m1_r1_cfg_1),
      .o_dq_dq_rx_io_m1_r1_cfg_2 (o_dq_dq_rx_io_m1_r1_cfg_2),
      .o_dq_dq_rx_io_m1_r1_cfg_3 (o_dq_dq_rx_io_m1_r1_cfg_3),
      .o_dq_dq_rx_io_m1_r1_cfg_4 (o_dq_dq_rx_io_m1_r1_cfg_4),
      .o_dq_dq_rx_io_m1_r1_cfg_5 (o_dq_dq_rx_io_m1_r1_cfg_5),
      .o_dq_dq_rx_io_m1_r1_cfg_6 (o_dq_dq_rx_io_m1_r1_cfg_6),
      .o_dq_dq_rx_io_m1_r1_cfg_7 (o_dq_dq_rx_io_m1_r1_cfg_7),
      .o_dq_dq_rx_io_m1_r1_cfg_8 (o_dq_dq_rx_io_m1_r1_cfg_8),
      .i_dq_dq_rx_io_sta (i_dq_dq_rx_io_sta),
      .o_dq_dq_rx_sa_m0_r0_cfg_0 (o_dq_dq_rx_sa_m0_r0_cfg_0),
      .o_dq_dq_rx_sa_m0_r0_cfg_1 (o_dq_dq_rx_sa_m0_r0_cfg_1),
      .o_dq_dq_rx_sa_m0_r0_cfg_2 (o_dq_dq_rx_sa_m0_r0_cfg_2),
      .o_dq_dq_rx_sa_m0_r0_cfg_3 (o_dq_dq_rx_sa_m0_r0_cfg_3),
      .o_dq_dq_rx_sa_m0_r0_cfg_4 (o_dq_dq_rx_sa_m0_r0_cfg_4),
      .o_dq_dq_rx_sa_m0_r0_cfg_5 (o_dq_dq_rx_sa_m0_r0_cfg_5),
      .o_dq_dq_rx_sa_m0_r0_cfg_6 (o_dq_dq_rx_sa_m0_r0_cfg_6),
      .o_dq_dq_rx_sa_m0_r0_cfg_7 (o_dq_dq_rx_sa_m0_r0_cfg_7),
      .o_dq_dq_rx_sa_m0_r0_cfg_8 (o_dq_dq_rx_sa_m0_r0_cfg_8),
      .o_dq_dq_rx_sa_m0_r1_cfg_0 (o_dq_dq_rx_sa_m0_r1_cfg_0),
      .o_dq_dq_rx_sa_m0_r1_cfg_1 (o_dq_dq_rx_sa_m0_r1_cfg_1),
      .o_dq_dq_rx_sa_m0_r1_cfg_2 (o_dq_dq_rx_sa_m0_r1_cfg_2),
      .o_dq_dq_rx_sa_m0_r1_cfg_3 (o_dq_dq_rx_sa_m0_r1_cfg_3),
      .o_dq_dq_rx_sa_m0_r1_cfg_4 (o_dq_dq_rx_sa_m0_r1_cfg_4),
      .o_dq_dq_rx_sa_m0_r1_cfg_5 (o_dq_dq_rx_sa_m0_r1_cfg_5),
      .o_dq_dq_rx_sa_m0_r1_cfg_6 (o_dq_dq_rx_sa_m0_r1_cfg_6),
      .o_dq_dq_rx_sa_m0_r1_cfg_7 (o_dq_dq_rx_sa_m0_r1_cfg_7),
      .o_dq_dq_rx_sa_m0_r1_cfg_8 (o_dq_dq_rx_sa_m0_r1_cfg_8),
      .o_dq_dq_rx_sa_m1_r0_cfg_0 (o_dq_dq_rx_sa_m1_r0_cfg_0),
      .o_dq_dq_rx_sa_m1_r0_cfg_1 (o_dq_dq_rx_sa_m1_r0_cfg_1),
      .o_dq_dq_rx_sa_m1_r0_cfg_2 (o_dq_dq_rx_sa_m1_r0_cfg_2),
      .o_dq_dq_rx_sa_m1_r0_cfg_3 (o_dq_dq_rx_sa_m1_r0_cfg_3),
      .o_dq_dq_rx_sa_m1_r0_cfg_4 (o_dq_dq_rx_sa_m1_r0_cfg_4),
      .o_dq_dq_rx_sa_m1_r0_cfg_5 (o_dq_dq_rx_sa_m1_r0_cfg_5),
      .o_dq_dq_rx_sa_m1_r0_cfg_6 (o_dq_dq_rx_sa_m1_r0_cfg_6),
      .o_dq_dq_rx_sa_m1_r0_cfg_7 (o_dq_dq_rx_sa_m1_r0_cfg_7),
      .o_dq_dq_rx_sa_m1_r0_cfg_8 (o_dq_dq_rx_sa_m1_r0_cfg_8),
      .o_dq_dq_rx_sa_m1_r1_cfg_0 (o_dq_dq_rx_sa_m1_r1_cfg_0),
      .o_dq_dq_rx_sa_m1_r1_cfg_1 (o_dq_dq_rx_sa_m1_r1_cfg_1),
      .o_dq_dq_rx_sa_m1_r1_cfg_2 (o_dq_dq_rx_sa_m1_r1_cfg_2),
      .o_dq_dq_rx_sa_m1_r1_cfg_3 (o_dq_dq_rx_sa_m1_r1_cfg_3),
      .o_dq_dq_rx_sa_m1_r1_cfg_4 (o_dq_dq_rx_sa_m1_r1_cfg_4),
      .o_dq_dq_rx_sa_m1_r1_cfg_5 (o_dq_dq_rx_sa_m1_r1_cfg_5),
      .o_dq_dq_rx_sa_m1_r1_cfg_6 (o_dq_dq_rx_sa_m1_r1_cfg_6),
      .o_dq_dq_rx_sa_m1_r1_cfg_7 (o_dq_dq_rx_sa_m1_r1_cfg_7),
      .o_dq_dq_rx_sa_m1_r1_cfg_8 (o_dq_dq_rx_sa_m1_r1_cfg_8),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_0 (o_dq_dq_rx_sa_dly_m0_r0_cfg_0),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_1 (o_dq_dq_rx_sa_dly_m0_r0_cfg_1),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_2 (o_dq_dq_rx_sa_dly_m0_r0_cfg_2),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_3 (o_dq_dq_rx_sa_dly_m0_r0_cfg_3),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_4 (o_dq_dq_rx_sa_dly_m0_r0_cfg_4),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_5 (o_dq_dq_rx_sa_dly_m0_r0_cfg_5),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_6 (o_dq_dq_rx_sa_dly_m0_r0_cfg_6),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_7 (o_dq_dq_rx_sa_dly_m0_r0_cfg_7),
      .o_dq_dq_rx_sa_dly_m0_r0_cfg_8 (o_dq_dq_rx_sa_dly_m0_r0_cfg_8),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_0 (o_dq_dq_rx_sa_dly_m0_r1_cfg_0),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_1 (o_dq_dq_rx_sa_dly_m0_r1_cfg_1),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_2 (o_dq_dq_rx_sa_dly_m0_r1_cfg_2),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_3 (o_dq_dq_rx_sa_dly_m0_r1_cfg_3),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_4 (o_dq_dq_rx_sa_dly_m0_r1_cfg_4),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_5 (o_dq_dq_rx_sa_dly_m0_r1_cfg_5),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_6 (o_dq_dq_rx_sa_dly_m0_r1_cfg_6),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_7 (o_dq_dq_rx_sa_dly_m0_r1_cfg_7),
      .o_dq_dq_rx_sa_dly_m0_r1_cfg_8 (o_dq_dq_rx_sa_dly_m0_r1_cfg_8),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_0 (o_dq_dq_rx_sa_dly_m1_r0_cfg_0),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_1 (o_dq_dq_rx_sa_dly_m1_r0_cfg_1),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_2 (o_dq_dq_rx_sa_dly_m1_r0_cfg_2),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_3 (o_dq_dq_rx_sa_dly_m1_r0_cfg_3),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_4 (o_dq_dq_rx_sa_dly_m1_r0_cfg_4),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_5 (o_dq_dq_rx_sa_dly_m1_r0_cfg_5),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_6 (o_dq_dq_rx_sa_dly_m1_r0_cfg_6),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_7 (o_dq_dq_rx_sa_dly_m1_r0_cfg_7),
      .o_dq_dq_rx_sa_dly_m1_r0_cfg_8 (o_dq_dq_rx_sa_dly_m1_r0_cfg_8),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_0 (o_dq_dq_rx_sa_dly_m1_r1_cfg_0),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_1 (o_dq_dq_rx_sa_dly_m1_r1_cfg_1),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_2 (o_dq_dq_rx_sa_dly_m1_r1_cfg_2),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_3 (o_dq_dq_rx_sa_dly_m1_r1_cfg_3),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_4 (o_dq_dq_rx_sa_dly_m1_r1_cfg_4),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_5 (o_dq_dq_rx_sa_dly_m1_r1_cfg_5),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_6 (o_dq_dq_rx_sa_dly_m1_r1_cfg_6),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_7 (o_dq_dq_rx_sa_dly_m1_r1_cfg_7),
      .o_dq_dq_rx_sa_dly_m1_r1_cfg_8 (o_dq_dq_rx_sa_dly_m1_r1_cfg_8),
      .i_dq_dq_rx_sa_sta_0 (i_dq_dq_rx_sa_sta_0),
      .i_dq_dq_rx_sa_sta_1 (i_dq_dq_rx_sa_sta_1),
      .i_dq_dq_rx_sa_sta_2 (i_dq_dq_rx_sa_sta_2),
      .i_dq_dq_rx_sa_sta_3 (i_dq_dq_rx_sa_sta_3),
      .i_dq_dq_rx_sa_sta_4 (i_dq_dq_rx_sa_sta_4),
      .i_dq_dq_rx_sa_sta_5 (i_dq_dq_rx_sa_sta_5),
      .i_dq_dq_rx_sa_sta_6 (i_dq_dq_rx_sa_sta_6),
      .i_dq_dq_rx_sa_sta_7 (i_dq_dq_rx_sa_sta_7),
      .i_dq_dq_rx_sa_sta_8 (i_dq_dq_rx_sa_sta_8),
      .o_dq_dq_tx_bscan_cfg (o_dq_dq_tx_bscan_cfg),
      .o_dq_dq_tx_egress_ana_m0_cfg_0 (o_dq_dq_tx_egress_ana_m0_cfg_0),
      .o_dq_dq_tx_egress_ana_m0_cfg_1 (o_dq_dq_tx_egress_ana_m0_cfg_1),
      .o_dq_dq_tx_egress_ana_m0_cfg_2 (o_dq_dq_tx_egress_ana_m0_cfg_2),
      .o_dq_dq_tx_egress_ana_m0_cfg_3 (o_dq_dq_tx_egress_ana_m0_cfg_3),
      .o_dq_dq_tx_egress_ana_m0_cfg_4 (o_dq_dq_tx_egress_ana_m0_cfg_4),
      .o_dq_dq_tx_egress_ana_m0_cfg_5 (o_dq_dq_tx_egress_ana_m0_cfg_5),
      .o_dq_dq_tx_egress_ana_m0_cfg_6 (o_dq_dq_tx_egress_ana_m0_cfg_6),
      .o_dq_dq_tx_egress_ana_m0_cfg_7 (o_dq_dq_tx_egress_ana_m0_cfg_7),
      .o_dq_dq_tx_egress_ana_m0_cfg_8 (o_dq_dq_tx_egress_ana_m0_cfg_8),
      .o_dq_dq_tx_egress_ana_m1_cfg_0 (o_dq_dq_tx_egress_ana_m1_cfg_0),
      .o_dq_dq_tx_egress_ana_m1_cfg_1 (o_dq_dq_tx_egress_ana_m1_cfg_1),
      .o_dq_dq_tx_egress_ana_m1_cfg_2 (o_dq_dq_tx_egress_ana_m1_cfg_2),
      .o_dq_dq_tx_egress_ana_m1_cfg_3 (o_dq_dq_tx_egress_ana_m1_cfg_3),
      .o_dq_dq_tx_egress_ana_m1_cfg_4 (o_dq_dq_tx_egress_ana_m1_cfg_4),
      .o_dq_dq_tx_egress_ana_m1_cfg_5 (o_dq_dq_tx_egress_ana_m1_cfg_5),
      .o_dq_dq_tx_egress_ana_m1_cfg_6 (o_dq_dq_tx_egress_ana_m1_cfg_6),
      .o_dq_dq_tx_egress_ana_m1_cfg_7 (o_dq_dq_tx_egress_ana_m1_cfg_7),
      .o_dq_dq_tx_egress_ana_m1_cfg_8 (o_dq_dq_tx_egress_ana_m1_cfg_8),
      .o_dq_dq_tx_egress_dig_m0_cfg_0 (o_dq_dq_tx_egress_dig_m0_cfg_0),
      .o_dq_dq_tx_egress_dig_m0_cfg_1 (o_dq_dq_tx_egress_dig_m0_cfg_1),
      .o_dq_dq_tx_egress_dig_m0_cfg_2 (o_dq_dq_tx_egress_dig_m0_cfg_2),
      .o_dq_dq_tx_egress_dig_m0_cfg_3 (o_dq_dq_tx_egress_dig_m0_cfg_3),
      .o_dq_dq_tx_egress_dig_m0_cfg_4 (o_dq_dq_tx_egress_dig_m0_cfg_4),
      .o_dq_dq_tx_egress_dig_m0_cfg_5 (o_dq_dq_tx_egress_dig_m0_cfg_5),
      .o_dq_dq_tx_egress_dig_m0_cfg_6 (o_dq_dq_tx_egress_dig_m0_cfg_6),
      .o_dq_dq_tx_egress_dig_m0_cfg_7 (o_dq_dq_tx_egress_dig_m0_cfg_7),
      .o_dq_dq_tx_egress_dig_m0_cfg_8 (o_dq_dq_tx_egress_dig_m0_cfg_8),
      .o_dq_dq_tx_egress_dig_m1_cfg_0 (o_dq_dq_tx_egress_dig_m1_cfg_0),
      .o_dq_dq_tx_egress_dig_m1_cfg_1 (o_dq_dq_tx_egress_dig_m1_cfg_1),
      .o_dq_dq_tx_egress_dig_m1_cfg_2 (o_dq_dq_tx_egress_dig_m1_cfg_2),
      .o_dq_dq_tx_egress_dig_m1_cfg_3 (o_dq_dq_tx_egress_dig_m1_cfg_3),
      .o_dq_dq_tx_egress_dig_m1_cfg_4 (o_dq_dq_tx_egress_dig_m1_cfg_4),
      .o_dq_dq_tx_egress_dig_m1_cfg_5 (o_dq_dq_tx_egress_dig_m1_cfg_5),
      .o_dq_dq_tx_egress_dig_m1_cfg_6 (o_dq_dq_tx_egress_dig_m1_cfg_6),
      .o_dq_dq_tx_egress_dig_m1_cfg_7 (o_dq_dq_tx_egress_dig_m1_cfg_7),
      .o_dq_dq_tx_egress_dig_m1_cfg_8 (o_dq_dq_tx_egress_dig_m1_cfg_8),
      .o_dq_dq_tx_odr_pi_m0_r0_cfg (o_dq_dq_tx_odr_pi_m0_r0_cfg),
      .o_dq_dq_tx_odr_pi_m0_r1_cfg (o_dq_dq_tx_odr_pi_m0_r1_cfg),
      .o_dq_dq_tx_odr_pi_m1_r0_cfg (o_dq_dq_tx_odr_pi_m1_r0_cfg),
      .o_dq_dq_tx_odr_pi_m1_r1_cfg (o_dq_dq_tx_odr_pi_m1_r1_cfg),
      .o_dq_dq_tx_qdr_pi_0_m0_r0_cfg (o_dq_dq_tx_qdr_pi_0_m0_r0_cfg),
      .o_dq_dq_tx_qdr_pi_0_m0_r1_cfg (o_dq_dq_tx_qdr_pi_0_m0_r1_cfg),
      .o_dq_dq_tx_qdr_pi_0_m1_r0_cfg (o_dq_dq_tx_qdr_pi_0_m1_r0_cfg),
      .o_dq_dq_tx_qdr_pi_0_m1_r1_cfg (o_dq_dq_tx_qdr_pi_0_m1_r1_cfg),
      .o_dq_dq_tx_qdr_pi_1_m0_r0_cfg (o_dq_dq_tx_qdr_pi_1_m0_r0_cfg),
      .o_dq_dq_tx_qdr_pi_1_m0_r1_cfg (o_dq_dq_tx_qdr_pi_1_m0_r1_cfg),
      .o_dq_dq_tx_qdr_pi_1_m1_r0_cfg (o_dq_dq_tx_qdr_pi_1_m1_r0_cfg),
      .o_dq_dq_tx_qdr_pi_1_m1_r1_cfg (o_dq_dq_tx_qdr_pi_1_m1_r1_cfg),
      .o_dq_dq_tx_ddr_pi_0_m0_r0_cfg (o_dq_dq_tx_ddr_pi_0_m0_r0_cfg),
      .o_dq_dq_tx_ddr_pi_0_m0_r1_cfg (o_dq_dq_tx_ddr_pi_0_m0_r1_cfg),
      .o_dq_dq_tx_ddr_pi_0_m1_r0_cfg (o_dq_dq_tx_ddr_pi_0_m1_r0_cfg),
      .o_dq_dq_tx_ddr_pi_0_m1_r1_cfg (o_dq_dq_tx_ddr_pi_0_m1_r1_cfg),
      .o_dq_dq_tx_ddr_pi_1_m0_r0_cfg (o_dq_dq_tx_ddr_pi_1_m0_r0_cfg),
      .o_dq_dq_tx_ddr_pi_1_m0_r1_cfg (o_dq_dq_tx_ddr_pi_1_m0_r1_cfg),
      .o_dq_dq_tx_ddr_pi_1_m1_r0_cfg (o_dq_dq_tx_ddr_pi_1_m1_r0_cfg),
      .o_dq_dq_tx_ddr_pi_1_m1_r1_cfg (o_dq_dq_tx_ddr_pi_1_m1_r1_cfg),
      .o_dq_dq_tx_pi_rt_m0_r0_cfg (o_dq_dq_tx_pi_rt_m0_r0_cfg),
      .o_dq_dq_tx_pi_rt_m0_r1_cfg (o_dq_dq_tx_pi_rt_m0_r1_cfg),
      .o_dq_dq_tx_pi_rt_m1_r0_cfg (o_dq_dq_tx_pi_rt_m1_r0_cfg),
      .o_dq_dq_tx_pi_rt_m1_r1_cfg (o_dq_dq_tx_pi_rt_m1_r1_cfg),
      .o_dq_dq_tx_rt_m0_r0_cfg (o_dq_dq_tx_rt_m0_r0_cfg),
      .o_dq_dq_tx_rt_m0_r1_cfg (o_dq_dq_tx_rt_m0_r1_cfg),
      .o_dq_dq_tx_rt_m1_r0_cfg (o_dq_dq_tx_rt_m1_r0_cfg),
      .o_dq_dq_tx_rt_m1_r1_cfg (o_dq_dq_tx_rt_m1_r1_cfg),
      .o_dq_dq_tx_sdr_m0_r0_cfg_0 (o_dq_dq_tx_sdr_m0_r0_cfg_0),
      .o_dq_dq_tx_sdr_m0_r0_cfg_1 (o_dq_dq_tx_sdr_m0_r0_cfg_1),
      .o_dq_dq_tx_sdr_m0_r0_cfg_2 (o_dq_dq_tx_sdr_m0_r0_cfg_2),
      .o_dq_dq_tx_sdr_m0_r0_cfg_3 (o_dq_dq_tx_sdr_m0_r0_cfg_3),
      .o_dq_dq_tx_sdr_m0_r0_cfg_4 (o_dq_dq_tx_sdr_m0_r0_cfg_4),
      .o_dq_dq_tx_sdr_m0_r0_cfg_5 (o_dq_dq_tx_sdr_m0_r0_cfg_5),
      .o_dq_dq_tx_sdr_m0_r0_cfg_6 (o_dq_dq_tx_sdr_m0_r0_cfg_6),
      .o_dq_dq_tx_sdr_m0_r0_cfg_7 (o_dq_dq_tx_sdr_m0_r0_cfg_7),
      .o_dq_dq_tx_sdr_m0_r0_cfg_8 (o_dq_dq_tx_sdr_m0_r0_cfg_8),
      .o_dq_dq_tx_sdr_m0_r1_cfg_0 (o_dq_dq_tx_sdr_m0_r1_cfg_0),
      .o_dq_dq_tx_sdr_m0_r1_cfg_1 (o_dq_dq_tx_sdr_m0_r1_cfg_1),
      .o_dq_dq_tx_sdr_m0_r1_cfg_2 (o_dq_dq_tx_sdr_m0_r1_cfg_2),
      .o_dq_dq_tx_sdr_m0_r1_cfg_3 (o_dq_dq_tx_sdr_m0_r1_cfg_3),
      .o_dq_dq_tx_sdr_m0_r1_cfg_4 (o_dq_dq_tx_sdr_m0_r1_cfg_4),
      .o_dq_dq_tx_sdr_m0_r1_cfg_5 (o_dq_dq_tx_sdr_m0_r1_cfg_5),
      .o_dq_dq_tx_sdr_m0_r1_cfg_6 (o_dq_dq_tx_sdr_m0_r1_cfg_6),
      .o_dq_dq_tx_sdr_m0_r1_cfg_7 (o_dq_dq_tx_sdr_m0_r1_cfg_7),
      .o_dq_dq_tx_sdr_m0_r1_cfg_8 (o_dq_dq_tx_sdr_m0_r1_cfg_8),
      .o_dq_dq_tx_sdr_m1_r0_cfg_0 (o_dq_dq_tx_sdr_m1_r0_cfg_0),
      .o_dq_dq_tx_sdr_m1_r0_cfg_1 (o_dq_dq_tx_sdr_m1_r0_cfg_1),
      .o_dq_dq_tx_sdr_m1_r0_cfg_2 (o_dq_dq_tx_sdr_m1_r0_cfg_2),
      .o_dq_dq_tx_sdr_m1_r0_cfg_3 (o_dq_dq_tx_sdr_m1_r0_cfg_3),
      .o_dq_dq_tx_sdr_m1_r0_cfg_4 (o_dq_dq_tx_sdr_m1_r0_cfg_4),
      .o_dq_dq_tx_sdr_m1_r0_cfg_5 (o_dq_dq_tx_sdr_m1_r0_cfg_5),
      .o_dq_dq_tx_sdr_m1_r0_cfg_6 (o_dq_dq_tx_sdr_m1_r0_cfg_6),
      .o_dq_dq_tx_sdr_m1_r0_cfg_7 (o_dq_dq_tx_sdr_m1_r0_cfg_7),
      .o_dq_dq_tx_sdr_m1_r0_cfg_8 (o_dq_dq_tx_sdr_m1_r0_cfg_8),
      .o_dq_dq_tx_sdr_m1_r1_cfg_0 (o_dq_dq_tx_sdr_m1_r1_cfg_0),
      .o_dq_dq_tx_sdr_m1_r1_cfg_1 (o_dq_dq_tx_sdr_m1_r1_cfg_1),
      .o_dq_dq_tx_sdr_m1_r1_cfg_2 (o_dq_dq_tx_sdr_m1_r1_cfg_2),
      .o_dq_dq_tx_sdr_m1_r1_cfg_3 (o_dq_dq_tx_sdr_m1_r1_cfg_3),
      .o_dq_dq_tx_sdr_m1_r1_cfg_4 (o_dq_dq_tx_sdr_m1_r1_cfg_4),
      .o_dq_dq_tx_sdr_m1_r1_cfg_5 (o_dq_dq_tx_sdr_m1_r1_cfg_5),
      .o_dq_dq_tx_sdr_m1_r1_cfg_6 (o_dq_dq_tx_sdr_m1_r1_cfg_6),
      .o_dq_dq_tx_sdr_m1_r1_cfg_7 (o_dq_dq_tx_sdr_m1_r1_cfg_7),
      .o_dq_dq_tx_sdr_m1_r1_cfg_8 (o_dq_dq_tx_sdr_m1_r1_cfg_8),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_0 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_0),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_1 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_1),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_2 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_2),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_3 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_3),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_4 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_4),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_5 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_5),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_6 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_6),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_7 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_7),
      .o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_8 (o_dq_dq_tx_sdr_x_sel_m0_r0_cfg_8),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_0 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_0),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_1 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_1),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_2 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_2),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_3 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_3),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_4 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_4),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_5 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_5),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_6 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_6),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_7 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_7),
      .o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_8 (o_dq_dq_tx_sdr_x_sel_m0_r1_cfg_8),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_0 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_0),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_1 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_1),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_2 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_2),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_3 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_3),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_4 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_4),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_5 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_5),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_6 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_6),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_7 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_7),
      .o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_8 (o_dq_dq_tx_sdr_x_sel_m1_r0_cfg_8),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_0 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_0),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_1 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_1),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_2 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_2),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_3 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_3),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_4 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_4),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_5 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_5),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_6 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_6),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_7 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_7),
      .o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_8 (o_dq_dq_tx_sdr_x_sel_m1_r1_cfg_8),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_0 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_0),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_1 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_1),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_2 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_2),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_3 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_3),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_4 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_4),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_5 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_5),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_6 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_6),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_7 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_7),
      .o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_8 (o_dq_dq_tx_sdr_fc_dly_m0_r0_cfg_8),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_0 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_0),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_1 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_1),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_2 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_2),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_3 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_3),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_4 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_4),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_5 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_5),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_6 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_6),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_7 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_7),
      .o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_8 (o_dq_dq_tx_sdr_fc_dly_m0_r1_cfg_8),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_0 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_0),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_1 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_1),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_2 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_2),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_3 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_3),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_4 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_4),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_5 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_5),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_6 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_6),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_7 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_7),
      .o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_8 (o_dq_dq_tx_sdr_fc_dly_m1_r0_cfg_8),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_0 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_0),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_1 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_1),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_2 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_2),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_3 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_3),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_4 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_4),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_5 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_5),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_6 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_6),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_7 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_7),
      .o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_8 (o_dq_dq_tx_sdr_fc_dly_m1_r1_cfg_8),
      .o_dq_dq_tx_ddr_m0_r0_cfg_0 (o_dq_dq_tx_ddr_m0_r0_cfg_0),
      .o_dq_dq_tx_ddr_m0_r0_cfg_1 (o_dq_dq_tx_ddr_m0_r0_cfg_1),
      .o_dq_dq_tx_ddr_m0_r0_cfg_2 (o_dq_dq_tx_ddr_m0_r0_cfg_2),
      .o_dq_dq_tx_ddr_m0_r0_cfg_3 (o_dq_dq_tx_ddr_m0_r0_cfg_3),
      .o_dq_dq_tx_ddr_m0_r0_cfg_4 (o_dq_dq_tx_ddr_m0_r0_cfg_4),
      .o_dq_dq_tx_ddr_m0_r0_cfg_5 (o_dq_dq_tx_ddr_m0_r0_cfg_5),
      .o_dq_dq_tx_ddr_m0_r0_cfg_6 (o_dq_dq_tx_ddr_m0_r0_cfg_6),
      .o_dq_dq_tx_ddr_m0_r0_cfg_7 (o_dq_dq_tx_ddr_m0_r0_cfg_7),
      .o_dq_dq_tx_ddr_m0_r0_cfg_8 (o_dq_dq_tx_ddr_m0_r0_cfg_8),
      .o_dq_dq_tx_ddr_m0_r1_cfg_0 (o_dq_dq_tx_ddr_m0_r1_cfg_0),
      .o_dq_dq_tx_ddr_m0_r1_cfg_1 (o_dq_dq_tx_ddr_m0_r1_cfg_1),
      .o_dq_dq_tx_ddr_m0_r1_cfg_2 (o_dq_dq_tx_ddr_m0_r1_cfg_2),
      .o_dq_dq_tx_ddr_m0_r1_cfg_3 (o_dq_dq_tx_ddr_m0_r1_cfg_3),
      .o_dq_dq_tx_ddr_m0_r1_cfg_4 (o_dq_dq_tx_ddr_m0_r1_cfg_4),
      .o_dq_dq_tx_ddr_m0_r1_cfg_5 (o_dq_dq_tx_ddr_m0_r1_cfg_5),
      .o_dq_dq_tx_ddr_m0_r1_cfg_6 (o_dq_dq_tx_ddr_m0_r1_cfg_6),
      .o_dq_dq_tx_ddr_m0_r1_cfg_7 (o_dq_dq_tx_ddr_m0_r1_cfg_7),
      .o_dq_dq_tx_ddr_m0_r1_cfg_8 (o_dq_dq_tx_ddr_m0_r1_cfg_8),
      .o_dq_dq_tx_ddr_m1_r0_cfg_0 (o_dq_dq_tx_ddr_m1_r0_cfg_0),
      .o_dq_dq_tx_ddr_m1_r0_cfg_1 (o_dq_dq_tx_ddr_m1_r0_cfg_1),
      .o_dq_dq_tx_ddr_m1_r0_cfg_2 (o_dq_dq_tx_ddr_m1_r0_cfg_2),
      .o_dq_dq_tx_ddr_m1_r0_cfg_3 (o_dq_dq_tx_ddr_m1_r0_cfg_3),
      .o_dq_dq_tx_ddr_m1_r0_cfg_4 (o_dq_dq_tx_ddr_m1_r0_cfg_4),
      .o_dq_dq_tx_ddr_m1_r0_cfg_5 (o_dq_dq_tx_ddr_m1_r0_cfg_5),
      .o_dq_dq_tx_ddr_m1_r0_cfg_6 (o_dq_dq_tx_ddr_m1_r0_cfg_6),
      .o_dq_dq_tx_ddr_m1_r0_cfg_7 (o_dq_dq_tx_ddr_m1_r0_cfg_7),
      .o_dq_dq_tx_ddr_m1_r0_cfg_8 (o_dq_dq_tx_ddr_m1_r0_cfg_8),
      .o_dq_dq_tx_ddr_m1_r1_cfg_0 (o_dq_dq_tx_ddr_m1_r1_cfg_0),
      .o_dq_dq_tx_ddr_m1_r1_cfg_1 (o_dq_dq_tx_ddr_m1_r1_cfg_1),
      .o_dq_dq_tx_ddr_m1_r1_cfg_2 (o_dq_dq_tx_ddr_m1_r1_cfg_2),
      .o_dq_dq_tx_ddr_m1_r1_cfg_3 (o_dq_dq_tx_ddr_m1_r1_cfg_3),
      .o_dq_dq_tx_ddr_m1_r1_cfg_4 (o_dq_dq_tx_ddr_m1_r1_cfg_4),
      .o_dq_dq_tx_ddr_m1_r1_cfg_5 (o_dq_dq_tx_ddr_m1_r1_cfg_5),
      .o_dq_dq_tx_ddr_m1_r1_cfg_6 (o_dq_dq_tx_ddr_m1_r1_cfg_6),
      .o_dq_dq_tx_ddr_m1_r1_cfg_7 (o_dq_dq_tx_ddr_m1_r1_cfg_7),
      .o_dq_dq_tx_ddr_m1_r1_cfg_8 (o_dq_dq_tx_ddr_m1_r1_cfg_8),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_0 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_0),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_1 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_1),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_2 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_2),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_3 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_3),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_4 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_4),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_5 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_5),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_6 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_6),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_7 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_7),
      .o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_8 (o_dq_dq_tx_ddr_x_sel_m0_r0_cfg_8),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_0 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_0),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_1 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_1),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_2 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_2),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_3 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_3),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_4 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_4),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_5 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_5),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_6 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_6),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_7 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_7),
      .o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_8 (o_dq_dq_tx_ddr_x_sel_m0_r1_cfg_8),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_0 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_0),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_1 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_1),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_2 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_2),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_3 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_3),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_4 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_4),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_5 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_5),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_6 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_6),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_7 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_7),
      .o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_8 (o_dq_dq_tx_ddr_x_sel_m1_r0_cfg_8),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_0 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_0),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_1 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_1),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_2 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_2),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_3 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_3),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_4 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_4),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_5 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_5),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_6 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_6),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_7 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_7),
      .o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_8 (o_dq_dq_tx_ddr_x_sel_m1_r1_cfg_8),
      .o_dq_dq_tx_qdr_m0_r0_cfg_0 (o_dq_dq_tx_qdr_m0_r0_cfg_0),
      .o_dq_dq_tx_qdr_m0_r0_cfg_1 (o_dq_dq_tx_qdr_m0_r0_cfg_1),
      .o_dq_dq_tx_qdr_m0_r0_cfg_2 (o_dq_dq_tx_qdr_m0_r0_cfg_2),
      .o_dq_dq_tx_qdr_m0_r0_cfg_3 (o_dq_dq_tx_qdr_m0_r0_cfg_3),
      .o_dq_dq_tx_qdr_m0_r0_cfg_4 (o_dq_dq_tx_qdr_m0_r0_cfg_4),
      .o_dq_dq_tx_qdr_m0_r0_cfg_5 (o_dq_dq_tx_qdr_m0_r0_cfg_5),
      .o_dq_dq_tx_qdr_m0_r0_cfg_6 (o_dq_dq_tx_qdr_m0_r0_cfg_6),
      .o_dq_dq_tx_qdr_m0_r0_cfg_7 (o_dq_dq_tx_qdr_m0_r0_cfg_7),
      .o_dq_dq_tx_qdr_m0_r0_cfg_8 (o_dq_dq_tx_qdr_m0_r0_cfg_8),
      .o_dq_dq_tx_qdr_m0_r1_cfg_0 (o_dq_dq_tx_qdr_m0_r1_cfg_0),
      .o_dq_dq_tx_qdr_m0_r1_cfg_1 (o_dq_dq_tx_qdr_m0_r1_cfg_1),
      .o_dq_dq_tx_qdr_m0_r1_cfg_2 (o_dq_dq_tx_qdr_m0_r1_cfg_2),
      .o_dq_dq_tx_qdr_m0_r1_cfg_3 (o_dq_dq_tx_qdr_m0_r1_cfg_3),
      .o_dq_dq_tx_qdr_m0_r1_cfg_4 (o_dq_dq_tx_qdr_m0_r1_cfg_4),
      .o_dq_dq_tx_qdr_m0_r1_cfg_5 (o_dq_dq_tx_qdr_m0_r1_cfg_5),
      .o_dq_dq_tx_qdr_m0_r1_cfg_6 (o_dq_dq_tx_qdr_m0_r1_cfg_6),
      .o_dq_dq_tx_qdr_m0_r1_cfg_7 (o_dq_dq_tx_qdr_m0_r1_cfg_7),
      .o_dq_dq_tx_qdr_m0_r1_cfg_8 (o_dq_dq_tx_qdr_m0_r1_cfg_8),
      .o_dq_dq_tx_qdr_m1_r0_cfg_0 (o_dq_dq_tx_qdr_m1_r0_cfg_0),
      .o_dq_dq_tx_qdr_m1_r0_cfg_1 (o_dq_dq_tx_qdr_m1_r0_cfg_1),
      .o_dq_dq_tx_qdr_m1_r0_cfg_2 (o_dq_dq_tx_qdr_m1_r0_cfg_2),
      .o_dq_dq_tx_qdr_m1_r0_cfg_3 (o_dq_dq_tx_qdr_m1_r0_cfg_3),
      .o_dq_dq_tx_qdr_m1_r0_cfg_4 (o_dq_dq_tx_qdr_m1_r0_cfg_4),
      .o_dq_dq_tx_qdr_m1_r0_cfg_5 (o_dq_dq_tx_qdr_m1_r0_cfg_5),
      .o_dq_dq_tx_qdr_m1_r0_cfg_6 (o_dq_dq_tx_qdr_m1_r0_cfg_6),
      .o_dq_dq_tx_qdr_m1_r0_cfg_7 (o_dq_dq_tx_qdr_m1_r0_cfg_7),
      .o_dq_dq_tx_qdr_m1_r0_cfg_8 (o_dq_dq_tx_qdr_m1_r0_cfg_8),
      .o_dq_dq_tx_qdr_m1_r1_cfg_0 (o_dq_dq_tx_qdr_m1_r1_cfg_0),
      .o_dq_dq_tx_qdr_m1_r1_cfg_1 (o_dq_dq_tx_qdr_m1_r1_cfg_1),
      .o_dq_dq_tx_qdr_m1_r1_cfg_2 (o_dq_dq_tx_qdr_m1_r1_cfg_2),
      .o_dq_dq_tx_qdr_m1_r1_cfg_3 (o_dq_dq_tx_qdr_m1_r1_cfg_3),
      .o_dq_dq_tx_qdr_m1_r1_cfg_4 (o_dq_dq_tx_qdr_m1_r1_cfg_4),
      .o_dq_dq_tx_qdr_m1_r1_cfg_5 (o_dq_dq_tx_qdr_m1_r1_cfg_5),
      .o_dq_dq_tx_qdr_m1_r1_cfg_6 (o_dq_dq_tx_qdr_m1_r1_cfg_6),
      .o_dq_dq_tx_qdr_m1_r1_cfg_7 (o_dq_dq_tx_qdr_m1_r1_cfg_7),
      .o_dq_dq_tx_qdr_m1_r1_cfg_8 (o_dq_dq_tx_qdr_m1_r1_cfg_8),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_0 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_0),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_1 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_1),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_2 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_2),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_3 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_3),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_4 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_4),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_5 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_5),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_6 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_6),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_7 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_7),
      .o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_8 (o_dq_dq_tx_qdr_x_sel_m0_r0_cfg_8),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_0 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_0),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_1 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_1),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_2 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_2),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_3 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_3),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_4 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_4),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_5 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_5),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_6 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_6),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_7 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_7),
      .o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_8 (o_dq_dq_tx_qdr_x_sel_m0_r1_cfg_8),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_0 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_0),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_1 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_1),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_2 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_2),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_3 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_3),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_4 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_4),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_5 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_5),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_6 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_6),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_7 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_7),
      .o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_8 (o_dq_dq_tx_qdr_x_sel_m1_r0_cfg_8),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_0 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_0),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_1 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_1),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_2 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_2),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_3 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_3),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_4 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_4),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_5 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_5),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_6 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_6),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_7 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_7),
      .o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_8 (o_dq_dq_tx_qdr_x_sel_m1_r1_cfg_8),
      .o_dq_dq_tx_lpde_m0_r0_cfg_0 (o_dq_dq_tx_lpde_m0_r0_cfg_0),
      .o_dq_dq_tx_lpde_m0_r0_cfg_1 (o_dq_dq_tx_lpde_m0_r0_cfg_1),
      .o_dq_dq_tx_lpde_m0_r0_cfg_2 (o_dq_dq_tx_lpde_m0_r0_cfg_2),
      .o_dq_dq_tx_lpde_m0_r0_cfg_3 (o_dq_dq_tx_lpde_m0_r0_cfg_3),
      .o_dq_dq_tx_lpde_m0_r0_cfg_4 (o_dq_dq_tx_lpde_m0_r0_cfg_4),
      .o_dq_dq_tx_lpde_m0_r0_cfg_5 (o_dq_dq_tx_lpde_m0_r0_cfg_5),
      .o_dq_dq_tx_lpde_m0_r0_cfg_6 (o_dq_dq_tx_lpde_m0_r0_cfg_6),
      .o_dq_dq_tx_lpde_m0_r0_cfg_7 (o_dq_dq_tx_lpde_m0_r0_cfg_7),
      .o_dq_dq_tx_lpde_m0_r0_cfg_8 (o_dq_dq_tx_lpde_m0_r0_cfg_8),
      .o_dq_dq_tx_lpde_m0_r1_cfg_0 (o_dq_dq_tx_lpde_m0_r1_cfg_0),
      .o_dq_dq_tx_lpde_m0_r1_cfg_1 (o_dq_dq_tx_lpde_m0_r1_cfg_1),
      .o_dq_dq_tx_lpde_m0_r1_cfg_2 (o_dq_dq_tx_lpde_m0_r1_cfg_2),
      .o_dq_dq_tx_lpde_m0_r1_cfg_3 (o_dq_dq_tx_lpde_m0_r1_cfg_3),
      .o_dq_dq_tx_lpde_m0_r1_cfg_4 (o_dq_dq_tx_lpde_m0_r1_cfg_4),
      .o_dq_dq_tx_lpde_m0_r1_cfg_5 (o_dq_dq_tx_lpde_m0_r1_cfg_5),
      .o_dq_dq_tx_lpde_m0_r1_cfg_6 (o_dq_dq_tx_lpde_m0_r1_cfg_6),
      .o_dq_dq_tx_lpde_m0_r1_cfg_7 (o_dq_dq_tx_lpde_m0_r1_cfg_7),
      .o_dq_dq_tx_lpde_m0_r1_cfg_8 (o_dq_dq_tx_lpde_m0_r1_cfg_8),
      .o_dq_dq_tx_lpde_m1_r0_cfg_0 (o_dq_dq_tx_lpde_m1_r0_cfg_0),
      .o_dq_dq_tx_lpde_m1_r0_cfg_1 (o_dq_dq_tx_lpde_m1_r0_cfg_1),
      .o_dq_dq_tx_lpde_m1_r0_cfg_2 (o_dq_dq_tx_lpde_m1_r0_cfg_2),
      .o_dq_dq_tx_lpde_m1_r0_cfg_3 (o_dq_dq_tx_lpde_m1_r0_cfg_3),
      .o_dq_dq_tx_lpde_m1_r0_cfg_4 (o_dq_dq_tx_lpde_m1_r0_cfg_4),
      .o_dq_dq_tx_lpde_m1_r0_cfg_5 (o_dq_dq_tx_lpde_m1_r0_cfg_5),
      .o_dq_dq_tx_lpde_m1_r0_cfg_6 (o_dq_dq_tx_lpde_m1_r0_cfg_6),
      .o_dq_dq_tx_lpde_m1_r0_cfg_7 (o_dq_dq_tx_lpde_m1_r0_cfg_7),
      .o_dq_dq_tx_lpde_m1_r0_cfg_8 (o_dq_dq_tx_lpde_m1_r0_cfg_8),
      .o_dq_dq_tx_lpde_m1_r1_cfg_0 (o_dq_dq_tx_lpde_m1_r1_cfg_0),
      .o_dq_dq_tx_lpde_m1_r1_cfg_1 (o_dq_dq_tx_lpde_m1_r1_cfg_1),
      .o_dq_dq_tx_lpde_m1_r1_cfg_2 (o_dq_dq_tx_lpde_m1_r1_cfg_2),
      .o_dq_dq_tx_lpde_m1_r1_cfg_3 (o_dq_dq_tx_lpde_m1_r1_cfg_3),
      .o_dq_dq_tx_lpde_m1_r1_cfg_4 (o_dq_dq_tx_lpde_m1_r1_cfg_4),
      .o_dq_dq_tx_lpde_m1_r1_cfg_5 (o_dq_dq_tx_lpde_m1_r1_cfg_5),
      .o_dq_dq_tx_lpde_m1_r1_cfg_6 (o_dq_dq_tx_lpde_m1_r1_cfg_6),
      .o_dq_dq_tx_lpde_m1_r1_cfg_7 (o_dq_dq_tx_lpde_m1_r1_cfg_7),
      .o_dq_dq_tx_lpde_m1_r1_cfg_8 (o_dq_dq_tx_lpde_m1_r1_cfg_8),
      .o_dq_dq_tx_io_m0_cfg_0 (o_dq_dq_tx_io_m0_cfg_0),
      .o_dq_dq_tx_io_m0_cfg_1 (o_dq_dq_tx_io_m0_cfg_1),
      .o_dq_dq_tx_io_m0_cfg_2 (o_dq_dq_tx_io_m0_cfg_2),
      .o_dq_dq_tx_io_m0_cfg_3 (o_dq_dq_tx_io_m0_cfg_3),
      .o_dq_dq_tx_io_m0_cfg_4 (o_dq_dq_tx_io_m0_cfg_4),
      .o_dq_dq_tx_io_m0_cfg_5 (o_dq_dq_tx_io_m0_cfg_5),
      .o_dq_dq_tx_io_m0_cfg_6 (o_dq_dq_tx_io_m0_cfg_6),
      .o_dq_dq_tx_io_m0_cfg_7 (o_dq_dq_tx_io_m0_cfg_7),
      .o_dq_dq_tx_io_m0_cfg_8 (o_dq_dq_tx_io_m0_cfg_8),
      .o_dq_dq_tx_io_m1_cfg_0 (o_dq_dq_tx_io_m1_cfg_0),
      .o_dq_dq_tx_io_m1_cfg_1 (o_dq_dq_tx_io_m1_cfg_1),
      .o_dq_dq_tx_io_m1_cfg_2 (o_dq_dq_tx_io_m1_cfg_2),
      .o_dq_dq_tx_io_m1_cfg_3 (o_dq_dq_tx_io_m1_cfg_3),
      .o_dq_dq_tx_io_m1_cfg_4 (o_dq_dq_tx_io_m1_cfg_4),
      .o_dq_dq_tx_io_m1_cfg_5 (o_dq_dq_tx_io_m1_cfg_5),
      .o_dq_dq_tx_io_m1_cfg_6 (o_dq_dq_tx_io_m1_cfg_6),
      .o_dq_dq_tx_io_m1_cfg_7 (o_dq_dq_tx_io_m1_cfg_7),
      .o_dq_dq_tx_io_m1_cfg_8 (o_dq_dq_tx_io_m1_cfg_8),
      .o_dq_dqs_rx_m0_cfg (o_dq_dqs_rx_m0_cfg),
      .o_dq_dqs_rx_m1_cfg (o_dq_dqs_rx_m1_cfg),
      .i_dq_dqs_rx_bscan_sta (i_dq_dqs_rx_bscan_sta),
      .o_dq_dqs_rx_sdr_lpde_m0_r0_cfg (o_dq_dqs_rx_sdr_lpde_m0_r0_cfg),
      .o_dq_dqs_rx_sdr_lpde_m0_r1_cfg (o_dq_dqs_rx_sdr_lpde_m0_r1_cfg),
      .o_dq_dqs_rx_sdr_lpde_m1_r0_cfg (o_dq_dqs_rx_sdr_lpde_m1_r0_cfg),
      .o_dq_dqs_rx_sdr_lpde_m1_r1_cfg (o_dq_dqs_rx_sdr_lpde_m1_r1_cfg),
      .o_dq_dqs_rx_ren_pi_m0_r0_cfg (o_dq_dqs_rx_ren_pi_m0_r0_cfg),
      .o_dq_dqs_rx_ren_pi_m0_r1_cfg (o_dq_dqs_rx_ren_pi_m0_r1_cfg),
      .o_dq_dqs_rx_ren_pi_m1_r0_cfg (o_dq_dqs_rx_ren_pi_m1_r0_cfg),
      .o_dq_dqs_rx_ren_pi_m1_r1_cfg (o_dq_dqs_rx_ren_pi_m1_r1_cfg),
      .o_dq_dqs_rx_rcs_pi_m0_r0_cfg (o_dq_dqs_rx_rcs_pi_m0_r0_cfg),
      .o_dq_dqs_rx_rcs_pi_m0_r1_cfg (o_dq_dqs_rx_rcs_pi_m0_r1_cfg),
      .o_dq_dqs_rx_rcs_pi_m1_r0_cfg (o_dq_dqs_rx_rcs_pi_m1_r0_cfg),
      .o_dq_dqs_rx_rcs_pi_m1_r1_cfg (o_dq_dqs_rx_rcs_pi_m1_r1_cfg),
      .o_dq_dqs_rx_rdqs_pi_0_m0_r0_cfg (o_dq_dqs_rx_rdqs_pi_0_m0_r0_cfg),
      .o_dq_dqs_rx_rdqs_pi_0_m0_r1_cfg (o_dq_dqs_rx_rdqs_pi_0_m0_r1_cfg),
      .o_dq_dqs_rx_rdqs_pi_0_m1_r0_cfg (o_dq_dqs_rx_rdqs_pi_0_m1_r0_cfg),
      .o_dq_dqs_rx_rdqs_pi_0_m1_r1_cfg (o_dq_dqs_rx_rdqs_pi_0_m1_r1_cfg),
      .o_dq_dqs_rx_rdqs_pi_1_m0_r0_cfg (o_dq_dqs_rx_rdqs_pi_1_m0_r0_cfg),
      .o_dq_dqs_rx_rdqs_pi_1_m0_r1_cfg (o_dq_dqs_rx_rdqs_pi_1_m0_r1_cfg),
      .o_dq_dqs_rx_rdqs_pi_1_m1_r0_cfg (o_dq_dqs_rx_rdqs_pi_1_m1_r0_cfg),
      .o_dq_dqs_rx_rdqs_pi_1_m1_r1_cfg (o_dq_dqs_rx_rdqs_pi_1_m1_r1_cfg),
      .i_dq_dqs_rx_pi_sta (i_dq_dqs_rx_pi_sta),
      .o_dq_dqs_rx_io_m0_r0_cfg_0 (o_dq_dqs_rx_io_m0_r0_cfg_0),
      .o_dq_dqs_rx_io_m0_r0_cfg_1 (o_dq_dqs_rx_io_m0_r0_cfg_1),
      .o_dq_dqs_rx_io_m0_r1_cfg_0 (o_dq_dqs_rx_io_m0_r1_cfg_0),
      .o_dq_dqs_rx_io_m0_r1_cfg_1 (o_dq_dqs_rx_io_m0_r1_cfg_1),
      .o_dq_dqs_rx_io_m1_r0_cfg_0 (o_dq_dqs_rx_io_m1_r0_cfg_0),
      .o_dq_dqs_rx_io_m1_r0_cfg_1 (o_dq_dqs_rx_io_m1_r0_cfg_1),
      .o_dq_dqs_rx_io_m1_r1_cfg_0 (o_dq_dqs_rx_io_m1_r1_cfg_0),
      .o_dq_dqs_rx_io_m1_r1_cfg_1 (o_dq_dqs_rx_io_m1_r1_cfg_1),
      .o_dq_dqs_rx_io_cmn_m0_r0_cfg (o_dq_dqs_rx_io_cmn_m0_r0_cfg),
      .o_dq_dqs_rx_io_cmn_m0_r1_cfg (o_dq_dqs_rx_io_cmn_m0_r1_cfg),
      .o_dq_dqs_rx_io_cmn_m1_r0_cfg (o_dq_dqs_rx_io_cmn_m1_r0_cfg),
      .o_dq_dqs_rx_io_cmn_m1_r1_cfg (o_dq_dqs_rx_io_cmn_m1_r1_cfg),
      .i_dq_dqs_rx_io_sta (i_dq_dqs_rx_io_sta),
      .o_dq_dqs_rx_sa_m0_r0_cfg_0 (o_dq_dqs_rx_sa_m0_r0_cfg_0),
      .o_dq_dqs_rx_sa_m0_r0_cfg_1 (o_dq_dqs_rx_sa_m0_r0_cfg_1),
      .o_dq_dqs_rx_sa_m0_r1_cfg_0 (o_dq_dqs_rx_sa_m0_r1_cfg_0),
      .o_dq_dqs_rx_sa_m0_r1_cfg_1 (o_dq_dqs_rx_sa_m0_r1_cfg_1),
      .o_dq_dqs_rx_sa_m1_r0_cfg_0 (o_dq_dqs_rx_sa_m1_r0_cfg_0),
      .o_dq_dqs_rx_sa_m1_r0_cfg_1 (o_dq_dqs_rx_sa_m1_r0_cfg_1),
      .o_dq_dqs_rx_sa_m1_r1_cfg_0 (o_dq_dqs_rx_sa_m1_r1_cfg_0),
      .o_dq_dqs_rx_sa_m1_r1_cfg_1 (o_dq_dqs_rx_sa_m1_r1_cfg_1),
      .o_dq_dqs_rx_sa_cmn_cfg (o_dq_dqs_rx_sa_cmn_cfg),
      .o_dq_dqs_tx_m0_cfg (o_dq_dqs_tx_m0_cfg),
      .o_dq_dqs_tx_m1_cfg (o_dq_dqs_tx_m1_cfg),
      .o_dq_dqs_tx_bscan_ctrl_cfg (o_dq_dqs_tx_bscan_ctrl_cfg),
      .o_dq_dqs_tx_bscan_cfg (o_dq_dqs_tx_bscan_cfg),
      .o_dq_dqs_tx_egress_ana_m0_cfg_0 (o_dq_dqs_tx_egress_ana_m0_cfg_0),
      .o_dq_dqs_tx_egress_ana_m0_cfg_1 (o_dq_dqs_tx_egress_ana_m0_cfg_1),
      .o_dq_dqs_tx_egress_ana_m0_cfg_2 (o_dq_dqs_tx_egress_ana_m0_cfg_2),
      .o_dq_dqs_tx_egress_ana_m0_cfg_3 (o_dq_dqs_tx_egress_ana_m0_cfg_3),
      .o_dq_dqs_tx_egress_ana_m0_cfg_4 (o_dq_dqs_tx_egress_ana_m0_cfg_4),
      .o_dq_dqs_tx_egress_ana_m0_cfg_5 (o_dq_dqs_tx_egress_ana_m0_cfg_5),
      .o_dq_dqs_tx_egress_ana_m0_cfg_6 (o_dq_dqs_tx_egress_ana_m0_cfg_6),
      .o_dq_dqs_tx_egress_ana_m0_cfg_7 (o_dq_dqs_tx_egress_ana_m0_cfg_7),
      .o_dq_dqs_tx_egress_ana_m0_cfg_8 (o_dq_dqs_tx_egress_ana_m0_cfg_8),
      .o_dq_dqs_tx_egress_ana_m1_cfg_0 (o_dq_dqs_tx_egress_ana_m1_cfg_0),
      .o_dq_dqs_tx_egress_ana_m1_cfg_1 (o_dq_dqs_tx_egress_ana_m1_cfg_1),
      .o_dq_dqs_tx_egress_ana_m1_cfg_2 (o_dq_dqs_tx_egress_ana_m1_cfg_2),
      .o_dq_dqs_tx_egress_ana_m1_cfg_3 (o_dq_dqs_tx_egress_ana_m1_cfg_3),
      .o_dq_dqs_tx_egress_ana_m1_cfg_4 (o_dq_dqs_tx_egress_ana_m1_cfg_4),
      .o_dq_dqs_tx_egress_ana_m1_cfg_5 (o_dq_dqs_tx_egress_ana_m1_cfg_5),
      .o_dq_dqs_tx_egress_ana_m1_cfg_6 (o_dq_dqs_tx_egress_ana_m1_cfg_6),
      .o_dq_dqs_tx_egress_ana_m1_cfg_7 (o_dq_dqs_tx_egress_ana_m1_cfg_7),
      .o_dq_dqs_tx_egress_ana_m1_cfg_8 (o_dq_dqs_tx_egress_ana_m1_cfg_8),
      .o_dq_dqs_tx_egress_dig_m0_cfg_0 (o_dq_dqs_tx_egress_dig_m0_cfg_0),
      .o_dq_dqs_tx_egress_dig_m0_cfg_1 (o_dq_dqs_tx_egress_dig_m0_cfg_1),
      .o_dq_dqs_tx_egress_dig_m0_cfg_2 (o_dq_dqs_tx_egress_dig_m0_cfg_2),
      .o_dq_dqs_tx_egress_dig_m0_cfg_3 (o_dq_dqs_tx_egress_dig_m0_cfg_3),
      .o_dq_dqs_tx_egress_dig_m0_cfg_4 (o_dq_dqs_tx_egress_dig_m0_cfg_4),
      .o_dq_dqs_tx_egress_dig_m0_cfg_5 (o_dq_dqs_tx_egress_dig_m0_cfg_5),
      .o_dq_dqs_tx_egress_dig_m0_cfg_6 (o_dq_dqs_tx_egress_dig_m0_cfg_6),
      .o_dq_dqs_tx_egress_dig_m0_cfg_7 (o_dq_dqs_tx_egress_dig_m0_cfg_7),
      .o_dq_dqs_tx_egress_dig_m0_cfg_8 (o_dq_dqs_tx_egress_dig_m0_cfg_8),
      .o_dq_dqs_tx_egress_dig_m1_cfg_0 (o_dq_dqs_tx_egress_dig_m1_cfg_0),
      .o_dq_dqs_tx_egress_dig_m1_cfg_1 (o_dq_dqs_tx_egress_dig_m1_cfg_1),
      .o_dq_dqs_tx_egress_dig_m1_cfg_2 (o_dq_dqs_tx_egress_dig_m1_cfg_2),
      .o_dq_dqs_tx_egress_dig_m1_cfg_3 (o_dq_dqs_tx_egress_dig_m1_cfg_3),
      .o_dq_dqs_tx_egress_dig_m1_cfg_4 (o_dq_dqs_tx_egress_dig_m1_cfg_4),
      .o_dq_dqs_tx_egress_dig_m1_cfg_5 (o_dq_dqs_tx_egress_dig_m1_cfg_5),
      .o_dq_dqs_tx_egress_dig_m1_cfg_6 (o_dq_dqs_tx_egress_dig_m1_cfg_6),
      .o_dq_dqs_tx_egress_dig_m1_cfg_7 (o_dq_dqs_tx_egress_dig_m1_cfg_7),
      .o_dq_dqs_tx_egress_dig_m1_cfg_8 (o_dq_dqs_tx_egress_dig_m1_cfg_8),
      .o_dq_dqs_tx_odr_pi_m0_r0_cfg (o_dq_dqs_tx_odr_pi_m0_r0_cfg),
      .o_dq_dqs_tx_odr_pi_m0_r1_cfg (o_dq_dqs_tx_odr_pi_m0_r1_cfg),
      .o_dq_dqs_tx_odr_pi_m1_r0_cfg (o_dq_dqs_tx_odr_pi_m1_r0_cfg),
      .o_dq_dqs_tx_odr_pi_m1_r1_cfg (o_dq_dqs_tx_odr_pi_m1_r1_cfg),
      .o_dq_dqs_tx_qdr_pi_0_m0_r0_cfg (o_dq_dqs_tx_qdr_pi_0_m0_r0_cfg),
      .o_dq_dqs_tx_qdr_pi_0_m0_r1_cfg (o_dq_dqs_tx_qdr_pi_0_m0_r1_cfg),
      .o_dq_dqs_tx_qdr_pi_0_m1_r0_cfg (o_dq_dqs_tx_qdr_pi_0_m1_r0_cfg),
      .o_dq_dqs_tx_qdr_pi_0_m1_r1_cfg (o_dq_dqs_tx_qdr_pi_0_m1_r1_cfg),
      .o_dq_dqs_tx_qdr_pi_1_m0_r0_cfg (o_dq_dqs_tx_qdr_pi_1_m0_r0_cfg),
      .o_dq_dqs_tx_qdr_pi_1_m0_r1_cfg (o_dq_dqs_tx_qdr_pi_1_m0_r1_cfg),
      .o_dq_dqs_tx_qdr_pi_1_m1_r0_cfg (o_dq_dqs_tx_qdr_pi_1_m1_r0_cfg),
      .o_dq_dqs_tx_qdr_pi_1_m1_r1_cfg (o_dq_dqs_tx_qdr_pi_1_m1_r1_cfg),
      .o_dq_dqs_tx_ddr_pi_0_m0_r0_cfg (o_dq_dqs_tx_ddr_pi_0_m0_r0_cfg),
      .o_dq_dqs_tx_ddr_pi_0_m0_r1_cfg (o_dq_dqs_tx_ddr_pi_0_m0_r1_cfg),
      .o_dq_dqs_tx_ddr_pi_0_m1_r0_cfg (o_dq_dqs_tx_ddr_pi_0_m1_r0_cfg),
      .o_dq_dqs_tx_ddr_pi_0_m1_r1_cfg (o_dq_dqs_tx_ddr_pi_0_m1_r1_cfg),
      .o_dq_dqs_tx_ddr_pi_1_m0_r0_cfg (o_dq_dqs_tx_ddr_pi_1_m0_r0_cfg),
      .o_dq_dqs_tx_ddr_pi_1_m0_r1_cfg (o_dq_dqs_tx_ddr_pi_1_m0_r1_cfg),
      .o_dq_dqs_tx_ddr_pi_1_m1_r0_cfg (o_dq_dqs_tx_ddr_pi_1_m1_r0_cfg),
      .o_dq_dqs_tx_ddr_pi_1_m1_r1_cfg (o_dq_dqs_tx_ddr_pi_1_m1_r1_cfg),
      .o_dq_dqs_tx_pi_rt_m0_r0_cfg (o_dq_dqs_tx_pi_rt_m0_r0_cfg),
      .o_dq_dqs_tx_pi_rt_m0_r1_cfg (o_dq_dqs_tx_pi_rt_m0_r1_cfg),
      .o_dq_dqs_tx_pi_rt_m1_r0_cfg (o_dq_dqs_tx_pi_rt_m1_r0_cfg),
      .o_dq_dqs_tx_pi_rt_m1_r1_cfg (o_dq_dqs_tx_pi_rt_m1_r1_cfg),
      .o_dq_dqs_tx_sdr_pi_m0_r0_cfg (o_dq_dqs_tx_sdr_pi_m0_r0_cfg),
      .o_dq_dqs_tx_sdr_pi_m0_r1_cfg (o_dq_dqs_tx_sdr_pi_m0_r1_cfg),
      .o_dq_dqs_tx_sdr_pi_m1_r0_cfg (o_dq_dqs_tx_sdr_pi_m1_r0_cfg),
      .o_dq_dqs_tx_sdr_pi_m1_r1_cfg (o_dq_dqs_tx_sdr_pi_m1_r1_cfg),
      .o_dq_dqs_tx_dfi_pi_m0_r0_cfg (o_dq_dqs_tx_dfi_pi_m0_r0_cfg),
      .o_dq_dqs_tx_dfi_pi_m0_r1_cfg (o_dq_dqs_tx_dfi_pi_m0_r1_cfg),
      .o_dq_dqs_tx_dfi_pi_m1_r0_cfg (o_dq_dqs_tx_dfi_pi_m1_r0_cfg),
      .o_dq_dqs_tx_dfi_pi_m1_r1_cfg (o_dq_dqs_tx_dfi_pi_m1_r1_cfg),
      .o_dq_dqs_tx_rt_m0_r0_cfg (o_dq_dqs_tx_rt_m0_r0_cfg),
      .o_dq_dqs_tx_rt_m0_r1_cfg (o_dq_dqs_tx_rt_m0_r1_cfg),
      .o_dq_dqs_tx_rt_m1_r0_cfg (o_dq_dqs_tx_rt_m1_r0_cfg),
      .o_dq_dqs_tx_rt_m1_r1_cfg (o_dq_dqs_tx_rt_m1_r1_cfg),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_0 (o_dq_dqs_tx_sdr_m0_r0_cfg_0),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_1 (o_dq_dqs_tx_sdr_m0_r0_cfg_1),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_2 (o_dq_dqs_tx_sdr_m0_r0_cfg_2),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_3 (o_dq_dqs_tx_sdr_m0_r0_cfg_3),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_4 (o_dq_dqs_tx_sdr_m0_r0_cfg_4),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_5 (o_dq_dqs_tx_sdr_m0_r0_cfg_5),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_6 (o_dq_dqs_tx_sdr_m0_r0_cfg_6),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_7 (o_dq_dqs_tx_sdr_m0_r0_cfg_7),
      .o_dq_dqs_tx_sdr_m0_r0_cfg_8 (o_dq_dqs_tx_sdr_m0_r0_cfg_8),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_0 (o_dq_dqs_tx_sdr_m0_r1_cfg_0),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_1 (o_dq_dqs_tx_sdr_m0_r1_cfg_1),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_2 (o_dq_dqs_tx_sdr_m0_r1_cfg_2),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_3 (o_dq_dqs_tx_sdr_m0_r1_cfg_3),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_4 (o_dq_dqs_tx_sdr_m0_r1_cfg_4),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_5 (o_dq_dqs_tx_sdr_m0_r1_cfg_5),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_6 (o_dq_dqs_tx_sdr_m0_r1_cfg_6),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_7 (o_dq_dqs_tx_sdr_m0_r1_cfg_7),
      .o_dq_dqs_tx_sdr_m0_r1_cfg_8 (o_dq_dqs_tx_sdr_m0_r1_cfg_8),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_0 (o_dq_dqs_tx_sdr_m1_r0_cfg_0),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_1 (o_dq_dqs_tx_sdr_m1_r0_cfg_1),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_2 (o_dq_dqs_tx_sdr_m1_r0_cfg_2),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_3 (o_dq_dqs_tx_sdr_m1_r0_cfg_3),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_4 (o_dq_dqs_tx_sdr_m1_r0_cfg_4),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_5 (o_dq_dqs_tx_sdr_m1_r0_cfg_5),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_6 (o_dq_dqs_tx_sdr_m1_r0_cfg_6),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_7 (o_dq_dqs_tx_sdr_m1_r0_cfg_7),
      .o_dq_dqs_tx_sdr_m1_r0_cfg_8 (o_dq_dqs_tx_sdr_m1_r0_cfg_8),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_0 (o_dq_dqs_tx_sdr_m1_r1_cfg_0),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_1 (o_dq_dqs_tx_sdr_m1_r1_cfg_1),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_2 (o_dq_dqs_tx_sdr_m1_r1_cfg_2),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_3 (o_dq_dqs_tx_sdr_m1_r1_cfg_3),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_4 (o_dq_dqs_tx_sdr_m1_r1_cfg_4),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_5 (o_dq_dqs_tx_sdr_m1_r1_cfg_5),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_6 (o_dq_dqs_tx_sdr_m1_r1_cfg_6),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_7 (o_dq_dqs_tx_sdr_m1_r1_cfg_7),
      .o_dq_dqs_tx_sdr_m1_r1_cfg_8 (o_dq_dqs_tx_sdr_m1_r1_cfg_8),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_0 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_0),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_1 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_1),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_2 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_2),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_3 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_3),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_4 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_4),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_5 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_5),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_6 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_6),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_7 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_7),
      .o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_8 (o_dq_dqs_tx_sdr_x_sel_m0_r0_cfg_8),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_0 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_0),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_1 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_1),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_2 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_2),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_3 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_3),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_4 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_4),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_5 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_5),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_6 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_6),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_7 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_7),
      .o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_8 (o_dq_dqs_tx_sdr_x_sel_m0_r1_cfg_8),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_0 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_0),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_1 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_1),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_2 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_2),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_3 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_3),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_4 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_4),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_5 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_5),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_6 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_6),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_7 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_7),
      .o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_8 (o_dq_dqs_tx_sdr_x_sel_m1_r0_cfg_8),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_0 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_0),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_1 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_1),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_2 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_2),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_3 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_3),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_4 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_4),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_5 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_5),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_6 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_6),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_7 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_7),
      .o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_8 (o_dq_dqs_tx_sdr_x_sel_m1_r1_cfg_8),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_0 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_0),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_1 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_1),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_2 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_2),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_3 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_3),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_4 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_4),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_5 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_5),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_6 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_6),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_7 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_7),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_8 (o_dq_dqs_tx_sdr_fc_dly_m0_r0_cfg_8),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_0 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_0),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_1 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_1),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_2 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_2),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_3 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_3),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_4 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_4),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_5 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_5),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_6 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_6),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_7 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_7),
      .o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_8 (o_dq_dqs_tx_sdr_fc_dly_m0_r1_cfg_8),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_0 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_0),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_1 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_1),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_2 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_2),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_3 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_3),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_4 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_4),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_5 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_5),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_6 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_6),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_7 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_7),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_8 (o_dq_dqs_tx_sdr_fc_dly_m1_r0_cfg_8),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_0 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_0),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_1 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_1),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_2 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_2),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_3 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_3),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_4 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_4),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_5 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_5),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_6 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_6),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_7 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_7),
      .o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_8 (o_dq_dqs_tx_sdr_fc_dly_m1_r1_cfg_8),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_0 (o_dq_dqs_tx_ddr_m0_r0_cfg_0),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_1 (o_dq_dqs_tx_ddr_m0_r0_cfg_1),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_2 (o_dq_dqs_tx_ddr_m0_r0_cfg_2),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_3 (o_dq_dqs_tx_ddr_m0_r0_cfg_3),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_4 (o_dq_dqs_tx_ddr_m0_r0_cfg_4),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_5 (o_dq_dqs_tx_ddr_m0_r0_cfg_5),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_6 (o_dq_dqs_tx_ddr_m0_r0_cfg_6),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_7 (o_dq_dqs_tx_ddr_m0_r0_cfg_7),
      .o_dq_dqs_tx_ddr_m0_r0_cfg_8 (o_dq_dqs_tx_ddr_m0_r0_cfg_8),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_0 (o_dq_dqs_tx_ddr_m0_r1_cfg_0),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_1 (o_dq_dqs_tx_ddr_m0_r1_cfg_1),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_2 (o_dq_dqs_tx_ddr_m0_r1_cfg_2),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_3 (o_dq_dqs_tx_ddr_m0_r1_cfg_3),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_4 (o_dq_dqs_tx_ddr_m0_r1_cfg_4),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_5 (o_dq_dqs_tx_ddr_m0_r1_cfg_5),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_6 (o_dq_dqs_tx_ddr_m0_r1_cfg_6),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_7 (o_dq_dqs_tx_ddr_m0_r1_cfg_7),
      .o_dq_dqs_tx_ddr_m0_r1_cfg_8 (o_dq_dqs_tx_ddr_m0_r1_cfg_8),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_0 (o_dq_dqs_tx_ddr_m1_r0_cfg_0),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_1 (o_dq_dqs_tx_ddr_m1_r0_cfg_1),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_2 (o_dq_dqs_tx_ddr_m1_r0_cfg_2),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_3 (o_dq_dqs_tx_ddr_m1_r0_cfg_3),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_4 (o_dq_dqs_tx_ddr_m1_r0_cfg_4),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_5 (o_dq_dqs_tx_ddr_m1_r0_cfg_5),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_6 (o_dq_dqs_tx_ddr_m1_r0_cfg_6),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_7 (o_dq_dqs_tx_ddr_m1_r0_cfg_7),
      .o_dq_dqs_tx_ddr_m1_r0_cfg_8 (o_dq_dqs_tx_ddr_m1_r0_cfg_8),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_0 (o_dq_dqs_tx_ddr_m1_r1_cfg_0),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_1 (o_dq_dqs_tx_ddr_m1_r1_cfg_1),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_2 (o_dq_dqs_tx_ddr_m1_r1_cfg_2),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_3 (o_dq_dqs_tx_ddr_m1_r1_cfg_3),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_4 (o_dq_dqs_tx_ddr_m1_r1_cfg_4),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_5 (o_dq_dqs_tx_ddr_m1_r1_cfg_5),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_6 (o_dq_dqs_tx_ddr_m1_r1_cfg_6),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_7 (o_dq_dqs_tx_ddr_m1_r1_cfg_7),
      .o_dq_dqs_tx_ddr_m1_r1_cfg_8 (o_dq_dqs_tx_ddr_m1_r1_cfg_8),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_0 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_0),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_1 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_1),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_2 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_2),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_3 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_3),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_4 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_4),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_5 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_5),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_6 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_6),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_7 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_7),
      .o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_8 (o_dq_dqs_tx_ddr_x_sel_m0_r0_cfg_8),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_0 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_0),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_1 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_1),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_2 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_2),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_3 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_3),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_4 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_4),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_5 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_5),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_6 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_6),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_7 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_7),
      .o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_8 (o_dq_dqs_tx_ddr_x_sel_m0_r1_cfg_8),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_0 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_0),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_1 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_1),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_2 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_2),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_3 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_3),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_4 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_4),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_5 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_5),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_6 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_6),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_7 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_7),
      .o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_8 (o_dq_dqs_tx_ddr_x_sel_m1_r0_cfg_8),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_0 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_0),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_1 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_1),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_2 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_2),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_3 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_3),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_4 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_4),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_5 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_5),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_6 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_6),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_7 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_7),
      .o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_8 (o_dq_dqs_tx_ddr_x_sel_m1_r1_cfg_8),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_0 (o_dq_dqs_tx_qdr_m0_r0_cfg_0),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_1 (o_dq_dqs_tx_qdr_m0_r0_cfg_1),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_2 (o_dq_dqs_tx_qdr_m0_r0_cfg_2),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_3 (o_dq_dqs_tx_qdr_m0_r0_cfg_3),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_4 (o_dq_dqs_tx_qdr_m0_r0_cfg_4),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_5 (o_dq_dqs_tx_qdr_m0_r0_cfg_5),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_6 (o_dq_dqs_tx_qdr_m0_r0_cfg_6),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_7 (o_dq_dqs_tx_qdr_m0_r0_cfg_7),
      .o_dq_dqs_tx_qdr_m0_r0_cfg_8 (o_dq_dqs_tx_qdr_m0_r0_cfg_8),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_0 (o_dq_dqs_tx_qdr_m0_r1_cfg_0),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_1 (o_dq_dqs_tx_qdr_m0_r1_cfg_1),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_2 (o_dq_dqs_tx_qdr_m0_r1_cfg_2),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_3 (o_dq_dqs_tx_qdr_m0_r1_cfg_3),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_4 (o_dq_dqs_tx_qdr_m0_r1_cfg_4),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_5 (o_dq_dqs_tx_qdr_m0_r1_cfg_5),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_6 (o_dq_dqs_tx_qdr_m0_r1_cfg_6),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_7 (o_dq_dqs_tx_qdr_m0_r1_cfg_7),
      .o_dq_dqs_tx_qdr_m0_r1_cfg_8 (o_dq_dqs_tx_qdr_m0_r1_cfg_8),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_0 (o_dq_dqs_tx_qdr_m1_r0_cfg_0),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_1 (o_dq_dqs_tx_qdr_m1_r0_cfg_1),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_2 (o_dq_dqs_tx_qdr_m1_r0_cfg_2),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_3 (o_dq_dqs_tx_qdr_m1_r0_cfg_3),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_4 (o_dq_dqs_tx_qdr_m1_r0_cfg_4),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_5 (o_dq_dqs_tx_qdr_m1_r0_cfg_5),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_6 (o_dq_dqs_tx_qdr_m1_r0_cfg_6),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_7 (o_dq_dqs_tx_qdr_m1_r0_cfg_7),
      .o_dq_dqs_tx_qdr_m1_r0_cfg_8 (o_dq_dqs_tx_qdr_m1_r0_cfg_8),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_0 (o_dq_dqs_tx_qdr_m1_r1_cfg_0),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_1 (o_dq_dqs_tx_qdr_m1_r1_cfg_1),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_2 (o_dq_dqs_tx_qdr_m1_r1_cfg_2),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_3 (o_dq_dqs_tx_qdr_m1_r1_cfg_3),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_4 (o_dq_dqs_tx_qdr_m1_r1_cfg_4),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_5 (o_dq_dqs_tx_qdr_m1_r1_cfg_5),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_6 (o_dq_dqs_tx_qdr_m1_r1_cfg_6),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_7 (o_dq_dqs_tx_qdr_m1_r1_cfg_7),
      .o_dq_dqs_tx_qdr_m1_r1_cfg_8 (o_dq_dqs_tx_qdr_m1_r1_cfg_8),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_0 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_0),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_1 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_1),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_2 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_2),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_3 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_3),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_4 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_4),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_5 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_5),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_6 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_6),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_7 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_7),
      .o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_8 (o_dq_dqs_tx_qdr_x_sel_m0_r0_cfg_8),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_0 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_0),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_1 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_1),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_2 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_2),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_3 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_3),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_4 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_4),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_5 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_5),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_6 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_6),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_7 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_7),
      .o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_8 (o_dq_dqs_tx_qdr_x_sel_m0_r1_cfg_8),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_0 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_0),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_1 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_1),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_2 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_2),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_3 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_3),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_4 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_4),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_5 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_5),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_6 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_6),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_7 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_7),
      .o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_8 (o_dq_dqs_tx_qdr_x_sel_m1_r0_cfg_8),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_0 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_0),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_1 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_1),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_2 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_2),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_3 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_3),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_4 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_4),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_5 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_5),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_6 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_6),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_7 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_7),
      .o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_8 (o_dq_dqs_tx_qdr_x_sel_m1_r1_cfg_8),
      .o_dq_dqs_tx_lpde_m0_r0_cfg_0 (o_dq_dqs_tx_lpde_m0_r0_cfg_0),
      .o_dq_dqs_tx_lpde_m0_r0_cfg_1 (o_dq_dqs_tx_lpde_m0_r0_cfg_1),
      .o_dq_dqs_tx_lpde_m0_r1_cfg_0 (o_dq_dqs_tx_lpde_m0_r1_cfg_0),
      .o_dq_dqs_tx_lpde_m0_r1_cfg_1 (o_dq_dqs_tx_lpde_m0_r1_cfg_1),
      .o_dq_dqs_tx_lpde_m1_r0_cfg_0 (o_dq_dqs_tx_lpde_m1_r0_cfg_0),
      .o_dq_dqs_tx_lpde_m1_r0_cfg_1 (o_dq_dqs_tx_lpde_m1_r0_cfg_1),
      .o_dq_dqs_tx_lpde_m1_r1_cfg_0 (o_dq_dqs_tx_lpde_m1_r1_cfg_0),
      .o_dq_dqs_tx_lpde_m1_r1_cfg_1 (o_dq_dqs_tx_lpde_m1_r1_cfg_1),
      .o_dq_dqs_tx_io_m0_cfg_0 (o_dq_dqs_tx_io_m0_cfg_0),
      .o_dq_dqs_tx_io_m0_cfg_1 (o_dq_dqs_tx_io_m0_cfg_1),
      .o_dq_dqs_tx_io_m1_cfg_0 (o_dq_dqs_tx_io_m1_cfg_0),
      .o_dq_dqs_tx_io_m1_cfg_1 (o_dq_dqs_tx_io_m1_cfg_1),
      .o_dq_dqs_tx_io_cmn_m0_r0_cfg (o_dq_dqs_tx_io_cmn_m0_r0_cfg),
      .o_dq_dqs_tx_io_cmn_m0_r1_cfg (o_dq_dqs_tx_io_cmn_m0_r1_cfg),
      .o_dq_dqs_tx_io_cmn_m1_r0_cfg (o_dq_dqs_tx_io_cmn_m1_r0_cfg),
      .o_dq_dqs_tx_io_cmn_m1_r1_cfg (o_dq_dqs_tx_io_cmn_m1_r1_cfg)
   );

endmodule
