/****************************************************************************
*****************************************************************************
** Wavious LLC Proprietary
**
** Copyright (c) 2019 Wavious LLC. All rights reserved.
**
** All data and information contained in or disclosed by this document
** are confidential and proprietary information of Wavious LLC,
** and all rights therein are expressly reserved. By accepting this
** material, the recipient agrees that this material and the information
** contained therein are held in confidence and in trust and will not be
** used, copied, reproduced in whole or in part, nor its contents
** revealed in any manner to others without the express written
** permission of Wavious LLC.
****************************************************************************
*
* Module    : ddr_ca_csr_defs.vh
* Date      : 2021-04-22
* Desciption: Autogenerated CSR block.
*
* $Id: ddr_ca_csr_defs.vh,v 1.109 2021/04/23 22:16:10 mclovis Exp $
*
****************************************************************************/

// Word Address 0x00000000 : DDR_CA_TOP_CFG (RW)
`define DDR_CA_TOP_CFG_FIFO_CLR_FIELD 8
`define DDR_CA_TOP_CFG_FIFO_CLR_FIELD_WIDTH 1
`define DDR_CA_TOP_CFG_RCS_SW_OVR_FIELD 2
`define DDR_CA_TOP_CFG_RCS_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_TOP_CFG_RCS_SW_OVR_VAL_FIELD 3
`define DDR_CA_TOP_CFG_RCS_SW_OVR_VAL_FIELD_WIDTH 1
`define DDR_CA_TOP_CFG_TRAINING_MODE_FIELD 9
`define DDR_CA_TOP_CFG_TRAINING_MODE_FIELD_WIDTH 1
`define DDR_CA_TOP_CFG_WCS_SW_OVR_FIELD 0
`define DDR_CA_TOP_CFG_WCS_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_TOP_CFG_WCS_SW_OVR_VAL_FIELD 1
`define DDR_CA_TOP_CFG_WCS_SW_OVR_VAL_FIELD_WIDTH 1
`define DDR_CA_TOP_CFG_RANGE 9:0
`define DDR_CA_TOP_CFG_WIDTH 10
`define DDR_CA_TOP_CFG_ADR 32'h00000000
`define DDR_CA_TOP_CFG_POR 32'h00000000
`define DDR_CA_TOP_CFG_MSK 32'h0000030F

// Word Address 0x00000004 : DDR_CA_TOP_STA (R)
`define DDR_CA_TOP_STA_RCS_FIELD 1
`define DDR_CA_TOP_STA_RCS_FIELD_WIDTH 1
`define DDR_CA_TOP_STA_WCS_FIELD 0
`define DDR_CA_TOP_STA_WCS_FIELD_WIDTH 1
`define DDR_CA_TOP_STA_RANGE 1:0
`define DDR_CA_TOP_STA_WIDTH 2
`define DDR_CA_TOP_STA_ADR 32'h00000004
`define DDR_CA_TOP_STA_POR 32'h00000000
`define DDR_CA_TOP_STA_MSK 32'h00000003

// Word Address 0x00000008 : DDR_CA_DQ_RX_BSCAN_STA (R)
`define DDR_CA_DQ_RX_BSCAN_STA_VAL_FIELD 10:0
`define DDR_CA_DQ_RX_BSCAN_STA_VAL_FIELD_WIDTH 11
`define DDR_CA_DQ_RX_BSCAN_STA_RANGE 10:0
`define DDR_CA_DQ_RX_BSCAN_STA_WIDTH 11
`define DDR_CA_DQ_RX_BSCAN_STA_ADR 32'h00000008
`define DDR_CA_DQ_RX_BSCAN_STA_POR 32'h00000000
`define DDR_CA_DQ_RX_BSCAN_STA_MSK 32'h000007FF

// Word Address 0x0000000C : DDR_CA_DQ_RX_M0_CFG (RW)
`define DDR_CA_DQ_RX_M0_CFG_FGB_MODE_FIELD 7:4
`define DDR_CA_DQ_RX_M0_CFG_FGB_MODE_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_M0_CFG_RGB_MODE_FIELD 2:0
`define DDR_CA_DQ_RX_M0_CFG_RGB_MODE_FIELD_WIDTH 3
`define DDR_CA_DQ_RX_M0_CFG_RANGE 7:0
`define DDR_CA_DQ_RX_M0_CFG_WIDTH 8
`define DDR_CA_DQ_RX_M0_CFG_ADR 32'h0000000C
`define DDR_CA_DQ_RX_M0_CFG_POR 32'h00000074
`define DDR_CA_DQ_RX_M0_CFG_MSK 32'h000000F7

// Word Address 0x00000010 : DDR_CA_DQ_RX_M1_CFG (RW)
`define DDR_CA_DQ_RX_M1_CFG_FGB_MODE_FIELD 7:4
`define DDR_CA_DQ_RX_M1_CFG_FGB_MODE_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_M1_CFG_RGB_MODE_FIELD 2:0
`define DDR_CA_DQ_RX_M1_CFG_RGB_MODE_FIELD_WIDTH 3
`define DDR_CA_DQ_RX_M1_CFG_RANGE 7:0
`define DDR_CA_DQ_RX_M1_CFG_WIDTH 8
`define DDR_CA_DQ_RX_M1_CFG_ADR 32'h00000010
`define DDR_CA_DQ_RX_M1_CFG_POR 32'h00000074
`define DDR_CA_DQ_RX_M1_CFG_MSK 32'h000000F7

// Word Address 0x00000014 : DDR_CA_DQ_RX_IO_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_ADR 32'h00000014
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_0_MSK 32'h000000FF

// Word Address 0x00000018 : DDR_CA_DQ_RX_IO_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_ADR 32'h00000018
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_1_MSK 32'h000000FF

// Word Address 0x0000001C : DDR_CA_DQ_RX_IO_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_ADR 32'h0000001C
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_2_MSK 32'h000000FF

// Word Address 0x00000020 : DDR_CA_DQ_RX_IO_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_ADR 32'h00000020
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_3_MSK 32'h000000FF

// Word Address 0x00000024 : DDR_CA_DQ_RX_IO_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_ADR 32'h00000024
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_4_MSK 32'h000000FF

// Word Address 0x00000028 : DDR_CA_DQ_RX_IO_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_ADR 32'h00000028
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_5_MSK 32'h000000FF

// Word Address 0x0000002C : DDR_CA_DQ_RX_IO_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_ADR 32'h0000002C
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_6_MSK 32'h000000FF

// Word Address 0x00000030 : DDR_CA_DQ_RX_IO_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_ADR 32'h00000030
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_7_MSK 32'h000000FF

// Word Address 0x00000034 : DDR_CA_DQ_RX_IO_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_ADR 32'h00000034
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_8_MSK 32'h000000FF

// Word Address 0x00000038 : DDR_CA_DQ_RX_IO_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_ADR 32'h00000038
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_9_MSK 32'h000000FF

// Word Address 0x0000003C : DDR_CA_DQ_RX_IO_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_ADR 32'h0000003C
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R0_CFG_10_MSK 32'h000000FF

// Word Address 0x00000040 : DDR_CA_DQ_RX_IO_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_ADR 32'h00000040
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_0_MSK 32'h000000FF

// Word Address 0x00000044 : DDR_CA_DQ_RX_IO_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_ADR 32'h00000044
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_1_MSK 32'h000000FF

// Word Address 0x00000048 : DDR_CA_DQ_RX_IO_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_ADR 32'h00000048
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_2_MSK 32'h000000FF

// Word Address 0x0000004C : DDR_CA_DQ_RX_IO_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_ADR 32'h0000004C
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_3_MSK 32'h000000FF

// Word Address 0x00000050 : DDR_CA_DQ_RX_IO_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_ADR 32'h00000050
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_4_MSK 32'h000000FF

// Word Address 0x00000054 : DDR_CA_DQ_RX_IO_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_ADR 32'h00000054
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_5_MSK 32'h000000FF

// Word Address 0x00000058 : DDR_CA_DQ_RX_IO_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_ADR 32'h00000058
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_6_MSK 32'h000000FF

// Word Address 0x0000005C : DDR_CA_DQ_RX_IO_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_ADR 32'h0000005C
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_7_MSK 32'h000000FF

// Word Address 0x00000060 : DDR_CA_DQ_RX_IO_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_ADR 32'h00000060
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_8_MSK 32'h000000FF

// Word Address 0x00000064 : DDR_CA_DQ_RX_IO_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_ADR 32'h00000064
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_9_MSK 32'h000000FF

// Word Address 0x00000068 : DDR_CA_DQ_RX_IO_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_WIDTH 8
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_ADR 32'h00000068
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M0_R1_CFG_10_MSK 32'h000000FF

// Word Address 0x0000006C : DDR_CA_DQ_RX_IO_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_ADR 32'h0000006C
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_0_MSK 32'h000000FF

// Word Address 0x00000070 : DDR_CA_DQ_RX_IO_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_ADR 32'h00000070
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_1_MSK 32'h000000FF

// Word Address 0x00000074 : DDR_CA_DQ_RX_IO_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_ADR 32'h00000074
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_2_MSK 32'h000000FF

// Word Address 0x00000078 : DDR_CA_DQ_RX_IO_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_ADR 32'h00000078
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_3_MSK 32'h000000FF

// Word Address 0x0000007C : DDR_CA_DQ_RX_IO_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_ADR 32'h0000007C
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_4_MSK 32'h000000FF

// Word Address 0x00000080 : DDR_CA_DQ_RX_IO_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_ADR 32'h00000080
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_5_MSK 32'h000000FF

// Word Address 0x00000084 : DDR_CA_DQ_RX_IO_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_ADR 32'h00000084
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_6_MSK 32'h000000FF

// Word Address 0x00000088 : DDR_CA_DQ_RX_IO_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_ADR 32'h00000088
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_7_MSK 32'h000000FF

// Word Address 0x0000008C : DDR_CA_DQ_RX_IO_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_ADR 32'h0000008C
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_8_MSK 32'h000000FF

// Word Address 0x00000090 : DDR_CA_DQ_RX_IO_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_ADR 32'h00000090
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_9_MSK 32'h000000FF

// Word Address 0x00000094 : DDR_CA_DQ_RX_IO_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_ADR 32'h00000094
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R0_CFG_10_MSK 32'h000000FF

// Word Address 0x00000098 : DDR_CA_DQ_RX_IO_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_ADR 32'h00000098
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_0_MSK 32'h000000FF

// Word Address 0x0000009C : DDR_CA_DQ_RX_IO_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_ADR 32'h0000009C
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_1_MSK 32'h000000FF

// Word Address 0x000000A0 : DDR_CA_DQ_RX_IO_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_ADR 32'h000000A0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_2_MSK 32'h000000FF

// Word Address 0x000000A4 : DDR_CA_DQ_RX_IO_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_ADR 32'h000000A4
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_3_MSK 32'h000000FF

// Word Address 0x000000A8 : DDR_CA_DQ_RX_IO_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_ADR 32'h000000A8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_4_MSK 32'h000000FF

// Word Address 0x000000AC : DDR_CA_DQ_RX_IO_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_ADR 32'h000000AC
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_5_MSK 32'h000000FF

// Word Address 0x000000B0 : DDR_CA_DQ_RX_IO_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_ADR 32'h000000B0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_6_MSK 32'h000000FF

// Word Address 0x000000B4 : DDR_CA_DQ_RX_IO_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_ADR 32'h000000B4
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_7_MSK 32'h000000FF

// Word Address 0x000000B8 : DDR_CA_DQ_RX_IO_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_ADR 32'h000000B8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_8_MSK 32'h000000FF

// Word Address 0x000000BC : DDR_CA_DQ_RX_IO_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_ADR 32'h000000BC
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_9_MSK 32'h000000FF

// Word Address 0x000000C0 : DDR_CA_DQ_RX_IO_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_RESERVED_FIELD 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_RESERVED_FIELD_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_RANGE 7:0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_WIDTH 8
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_ADR 32'h000000C0
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_M1_R1_CFG_10_MSK 32'h000000FF

// Word Address 0x000000C4 : DDR_CA_DQ_RX_IO_STA (R)
`define DDR_CA_DQ_RX_IO_STA_CORE_IG_FIELD 31:0
`define DDR_CA_DQ_RX_IO_STA_CORE_IG_FIELD_WIDTH 32
`define DDR_CA_DQ_RX_IO_STA_RANGE 31:0
`define DDR_CA_DQ_RX_IO_STA_WIDTH 32
`define DDR_CA_DQ_RX_IO_STA_ADR 32'h000000C4
`define DDR_CA_DQ_RX_IO_STA_POR 32'h00000000
`define DDR_CA_DQ_RX_IO_STA_MSK 32'hFFFFFFFF

// Word Address 0x000000C8 : DDR_CA_DQ_RX_SA_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_ADR 32'h000000C8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_0_MSK 32'h000FFFFF

// Word Address 0x000000CC : DDR_CA_DQ_RX_SA_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_ADR 32'h000000CC
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_1_MSK 32'h000FFFFF

// Word Address 0x000000D0 : DDR_CA_DQ_RX_SA_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_ADR 32'h000000D0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_2_MSK 32'h000FFFFF

// Word Address 0x000000D4 : DDR_CA_DQ_RX_SA_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_ADR 32'h000000D4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_3_MSK 32'h000FFFFF

// Word Address 0x000000D8 : DDR_CA_DQ_RX_SA_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_ADR 32'h000000D8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_4_MSK 32'h000FFFFF

// Word Address 0x000000DC : DDR_CA_DQ_RX_SA_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_ADR 32'h000000DC
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_5_MSK 32'h000FFFFF

// Word Address 0x000000E0 : DDR_CA_DQ_RX_SA_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_ADR 32'h000000E0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_6_MSK 32'h000FFFFF

// Word Address 0x000000E4 : DDR_CA_DQ_RX_SA_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_ADR 32'h000000E4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_7_MSK 32'h000FFFFF

// Word Address 0x000000E8 : DDR_CA_DQ_RX_SA_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_ADR 32'h000000E8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_8_MSK 32'h000FFFFF

// Word Address 0x000000EC : DDR_CA_DQ_RX_SA_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_ADR 32'h000000EC
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_9_MSK 32'h000FFFFF

// Word Address 0x000000F0 : DDR_CA_DQ_RX_SA_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_ADR 32'h000000F0
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R0_CFG_10_MSK 32'h000FFFFF

// Word Address 0x000000F4 : DDR_CA_DQ_RX_SA_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_ADR 32'h000000F4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_0_MSK 32'h000FFFFF

// Word Address 0x000000F8 : DDR_CA_DQ_RX_SA_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_ADR 32'h000000F8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_1_MSK 32'h000FFFFF

// Word Address 0x000000FC : DDR_CA_DQ_RX_SA_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_ADR 32'h000000FC
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_2_MSK 32'h000FFFFF

// Word Address 0x00000100 : DDR_CA_DQ_RX_SA_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_ADR 32'h00000100
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_3_MSK 32'h000FFFFF

// Word Address 0x00000104 : DDR_CA_DQ_RX_SA_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_ADR 32'h00000104
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_4_MSK 32'h000FFFFF

// Word Address 0x00000108 : DDR_CA_DQ_RX_SA_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_ADR 32'h00000108
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_5_MSK 32'h000FFFFF

// Word Address 0x0000010C : DDR_CA_DQ_RX_SA_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_ADR 32'h0000010C
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_6_MSK 32'h000FFFFF

// Word Address 0x00000110 : DDR_CA_DQ_RX_SA_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_ADR 32'h00000110
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_7_MSK 32'h000FFFFF

// Word Address 0x00000114 : DDR_CA_DQ_RX_SA_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_ADR 32'h00000114
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_8_MSK 32'h000FFFFF

// Word Address 0x00000118 : DDR_CA_DQ_RX_SA_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_ADR 32'h00000118
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_9_MSK 32'h000FFFFF

// Word Address 0x0000011C : DDR_CA_DQ_RX_SA_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_WIDTH 20
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_ADR 32'h0000011C
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M0_R1_CFG_10_MSK 32'h000FFFFF

// Word Address 0x00000120 : DDR_CA_DQ_RX_SA_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_ADR 32'h00000120
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_0_MSK 32'h000FFFFF

// Word Address 0x00000124 : DDR_CA_DQ_RX_SA_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_ADR 32'h00000124
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_1_MSK 32'h000FFFFF

// Word Address 0x00000128 : DDR_CA_DQ_RX_SA_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_ADR 32'h00000128
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_2_MSK 32'h000FFFFF

// Word Address 0x0000012C : DDR_CA_DQ_RX_SA_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_ADR 32'h0000012C
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_3_MSK 32'h000FFFFF

// Word Address 0x00000130 : DDR_CA_DQ_RX_SA_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_ADR 32'h00000130
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_4_MSK 32'h000FFFFF

// Word Address 0x00000134 : DDR_CA_DQ_RX_SA_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_ADR 32'h00000134
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_5_MSK 32'h000FFFFF

// Word Address 0x00000138 : DDR_CA_DQ_RX_SA_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_ADR 32'h00000138
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_6_MSK 32'h000FFFFF

// Word Address 0x0000013C : DDR_CA_DQ_RX_SA_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_ADR 32'h0000013C
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_7_MSK 32'h000FFFFF

// Word Address 0x00000140 : DDR_CA_DQ_RX_SA_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_ADR 32'h00000140
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_8_MSK 32'h000FFFFF

// Word Address 0x00000144 : DDR_CA_DQ_RX_SA_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_ADR 32'h00000144
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_9_MSK 32'h000FFFFF

// Word Address 0x00000148 : DDR_CA_DQ_RX_SA_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_ADR 32'h00000148
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R0_CFG_10_MSK 32'h000FFFFF

// Word Address 0x0000014C : DDR_CA_DQ_RX_SA_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_ADR 32'h0000014C
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_0_MSK 32'h000FFFFF

// Word Address 0x00000150 : DDR_CA_DQ_RX_SA_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_ADR 32'h00000150
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_1_MSK 32'h000FFFFF

// Word Address 0x00000154 : DDR_CA_DQ_RX_SA_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_ADR 32'h00000154
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_2_MSK 32'h000FFFFF

// Word Address 0x00000158 : DDR_CA_DQ_RX_SA_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_ADR 32'h00000158
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_3_MSK 32'h000FFFFF

// Word Address 0x0000015C : DDR_CA_DQ_RX_SA_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_ADR 32'h0000015C
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_4_MSK 32'h000FFFFF

// Word Address 0x00000160 : DDR_CA_DQ_RX_SA_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_ADR 32'h00000160
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_5_MSK 32'h000FFFFF

// Word Address 0x00000164 : DDR_CA_DQ_RX_SA_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_ADR 32'h00000164
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_6_MSK 32'h000FFFFF

// Word Address 0x00000168 : DDR_CA_DQ_RX_SA_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_ADR 32'h00000168
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_7_MSK 32'h000FFFFF

// Word Address 0x0000016C : DDR_CA_DQ_RX_SA_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_ADR 32'h0000016C
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_8_MSK 32'h000FFFFF

// Word Address 0x00000170 : DDR_CA_DQ_RX_SA_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_ADR 32'h00000170
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_9_MSK 32'h000FFFFF

// Word Address 0x00000174 : DDR_CA_DQ_RX_SA_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_0_FIELD 16
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_180_FIELD 18
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_270_FIELD 19
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_90_FIELD 17
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_RANGE 19:0
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_WIDTH 20
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_ADR 32'h00000174
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_M1_R1_CFG_10_MSK 32'h000FFFFF

// Word Address 0x00000178 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_ADR 32'h00000178
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_0_MSK 32'hFFFFFFFF

// Word Address 0x0000017C : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_ADR 32'h0000017C
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_1_MSK 32'hFFFFFFFF

// Word Address 0x00000180 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_ADR 32'h00000180
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_2_MSK 32'hFFFFFFFF

// Word Address 0x00000184 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_ADR 32'h00000184
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_3_MSK 32'hFFFFFFFF

// Word Address 0x00000188 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_ADR 32'h00000188
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_4_MSK 32'hFFFFFFFF

// Word Address 0x0000018C : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_ADR 32'h0000018C
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_5_MSK 32'hFFFFFFFF

// Word Address 0x00000190 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_ADR 32'h00000190
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_6_MSK 32'hFFFFFFFF

// Word Address 0x00000194 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_ADR 32'h00000194
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_7_MSK 32'hFFFFFFFF

// Word Address 0x00000198 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_ADR 32'h00000198
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_8_MSK 32'hFFFFFFFF

// Word Address 0x0000019C : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_ADR 32'h0000019C
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_9_MSK 32'hFFFFFFFF

// Word Address 0x000001A0 : DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_ADR 32'h000001A0
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R0_CFG_10_MSK 32'hFFFFFFFF

// Word Address 0x000001A4 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_ADR 32'h000001A4
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_0_MSK 32'hFFFFFFFF

// Word Address 0x000001A8 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_ADR 32'h000001A8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_1_MSK 32'hFFFFFFFF

// Word Address 0x000001AC : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_ADR 32'h000001AC
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_2_MSK 32'hFFFFFFFF

// Word Address 0x000001B0 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_ADR 32'h000001B0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_3_MSK 32'hFFFFFFFF

// Word Address 0x000001B4 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_ADR 32'h000001B4
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_4_MSK 32'hFFFFFFFF

// Word Address 0x000001B8 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_ADR 32'h000001B8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_5_MSK 32'hFFFFFFFF

// Word Address 0x000001BC : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_ADR 32'h000001BC
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_6_MSK 32'hFFFFFFFF

// Word Address 0x000001C0 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_ADR 32'h000001C0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_7_MSK 32'hFFFFFFFF

// Word Address 0x000001C4 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_ADR 32'h000001C4
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_8_MSK 32'hFFFFFFFF

// Word Address 0x000001C8 : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_ADR 32'h000001C8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_9_MSK 32'hFFFFFFFF

// Word Address 0x000001CC : DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_ADR 32'h000001CC
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M0_R1_CFG_10_MSK 32'hFFFFFFFF

// Word Address 0x000001D0 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_ADR 32'h000001D0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_0_MSK 32'hFFFFFFFF

// Word Address 0x000001D4 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_ADR 32'h000001D4
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_1_MSK 32'hFFFFFFFF

// Word Address 0x000001D8 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_ADR 32'h000001D8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_2_MSK 32'hFFFFFFFF

// Word Address 0x000001DC : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_ADR 32'h000001DC
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_3_MSK 32'hFFFFFFFF

// Word Address 0x000001E0 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_ADR 32'h000001E0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_4_MSK 32'hFFFFFFFF

// Word Address 0x000001E4 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_ADR 32'h000001E4
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_5_MSK 32'hFFFFFFFF

// Word Address 0x000001E8 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_ADR 32'h000001E8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_6_MSK 32'hFFFFFFFF

// Word Address 0x000001EC : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_ADR 32'h000001EC
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_7_MSK 32'hFFFFFFFF

// Word Address 0x000001F0 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_ADR 32'h000001F0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_8_MSK 32'hFFFFFFFF

// Word Address 0x000001F4 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_ADR 32'h000001F4
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_9_MSK 32'hFFFFFFFF

// Word Address 0x000001F8 : DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_ADR 32'h000001F8
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R0_CFG_10_MSK 32'hFFFFFFFF

// Word Address 0x000001FC : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_ADR 32'h000001FC
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_0_MSK 32'hFFFFFFFF

// Word Address 0x00000200 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_ADR 32'h00000200
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_1_MSK 32'hFFFFFFFF

// Word Address 0x00000204 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_ADR 32'h00000204
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_2_MSK 32'hFFFFFFFF

// Word Address 0x00000208 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_ADR 32'h00000208
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_3_MSK 32'hFFFFFFFF

// Word Address 0x0000020C : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_ADR 32'h0000020C
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_4_MSK 32'hFFFFFFFF

// Word Address 0x00000210 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_ADR 32'h00000210
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_5_MSK 32'hFFFFFFFF

// Word Address 0x00000214 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_ADR 32'h00000214
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_6_MSK 32'hFFFFFFFF

// Word Address 0x00000218 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_ADR 32'h00000218
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_7_MSK 32'hFFFFFFFF

// Word Address 0x0000021C : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_ADR 32'h0000021C
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_8_MSK 32'hFFFFFFFF

// Word Address 0x00000220 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_ADR 32'h00000220
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_9_MSK 32'hFFFFFFFF

// Word Address 0x00000224 : DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_0_FIELD 7:2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_0_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_180_FIELD 23:18
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_180_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_270_FIELD 31:26
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_270_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_90_FIELD 15:10
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_CTRL_90_FIELD_WIDTH 6
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_0_FIELD 1:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_0_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_180_FIELD 17:16
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_180_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_270_FIELD 25:24
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_270_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_90_FIELD 9:8
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_GEAR_90_FIELD_WIDTH 2
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_RANGE 31:0
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_WIDTH 32
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_ADR 32'h00000224
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_DLY_M1_R1_CFG_10_MSK 32'hFFFFFFFF

// Word Address 0x00000228 : DDR_CA_DQ_RX_SA_STA_0 (R)
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_0_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_0_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_0_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_0_ADR 32'h00000228
`define DDR_CA_DQ_RX_SA_STA_0_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_0_MSK 32'h0000000F

// Word Address 0x0000022C : DDR_CA_DQ_RX_SA_STA_1 (R)
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_1_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_1_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_1_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_1_ADR 32'h0000022C
`define DDR_CA_DQ_RX_SA_STA_1_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_1_MSK 32'h0000000F

// Word Address 0x00000230 : DDR_CA_DQ_RX_SA_STA_2 (R)
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_2_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_2_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_2_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_2_ADR 32'h00000230
`define DDR_CA_DQ_RX_SA_STA_2_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_2_MSK 32'h0000000F

// Word Address 0x00000234 : DDR_CA_DQ_RX_SA_STA_3 (R)
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_3_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_3_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_3_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_3_ADR 32'h00000234
`define DDR_CA_DQ_RX_SA_STA_3_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_3_MSK 32'h0000000F

// Word Address 0x00000238 : DDR_CA_DQ_RX_SA_STA_4 (R)
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_4_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_4_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_4_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_4_ADR 32'h00000238
`define DDR_CA_DQ_RX_SA_STA_4_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_4_MSK 32'h0000000F

// Word Address 0x0000023C : DDR_CA_DQ_RX_SA_STA_5 (R)
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_5_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_5_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_5_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_5_ADR 32'h0000023C
`define DDR_CA_DQ_RX_SA_STA_5_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_5_MSK 32'h0000000F

// Word Address 0x00000240 : DDR_CA_DQ_RX_SA_STA_6 (R)
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_6_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_6_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_6_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_6_ADR 32'h00000240
`define DDR_CA_DQ_RX_SA_STA_6_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_6_MSK 32'h0000000F

// Word Address 0x00000244 : DDR_CA_DQ_RX_SA_STA_7 (R)
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_7_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_7_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_7_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_7_ADR 32'h00000244
`define DDR_CA_DQ_RX_SA_STA_7_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_7_MSK 32'h0000000F

// Word Address 0x00000248 : DDR_CA_DQ_RX_SA_STA_8 (R)
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_8_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_8_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_8_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_8_ADR 32'h00000248
`define DDR_CA_DQ_RX_SA_STA_8_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_8_MSK 32'h0000000F

// Word Address 0x0000024C : DDR_CA_DQ_RX_SA_STA_9 (R)
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_9_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_9_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_9_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_9_ADR 32'h0000024C
`define DDR_CA_DQ_RX_SA_STA_9_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_9_MSK 32'h0000000F

// Word Address 0x00000250 : DDR_CA_DQ_RX_SA_STA_10 (R)
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_0_FIELD 0
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_0_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_180_FIELD 2
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_180_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_270_FIELD 3
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_270_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_90_FIELD 1
`define DDR_CA_DQ_RX_SA_STA_10_SA_OUT_90_FIELD_WIDTH 1
`define DDR_CA_DQ_RX_SA_STA_10_RANGE 3:0
`define DDR_CA_DQ_RX_SA_STA_10_WIDTH 4
`define DDR_CA_DQ_RX_SA_STA_10_ADR 32'h00000250
`define DDR_CA_DQ_RX_SA_STA_10_POR 32'h00000000
`define DDR_CA_DQ_RX_SA_STA_10_MSK 32'h0000000F

// Word Address 0x00000254 : DDR_CA_DQ_TX_BSCAN_CFG (RW)
`define DDR_CA_DQ_TX_BSCAN_CFG_VAL_FIELD 10:0
`define DDR_CA_DQ_TX_BSCAN_CFG_VAL_FIELD_WIDTH 11
`define DDR_CA_DQ_TX_BSCAN_CFG_RANGE 10:0
`define DDR_CA_DQ_TX_BSCAN_CFG_WIDTH 11
`define DDR_CA_DQ_TX_BSCAN_CFG_ADR 32'h00000254
`define DDR_CA_DQ_TX_BSCAN_CFG_POR 32'h00000000
`define DDR_CA_DQ_TX_BSCAN_CFG_MSK 32'h000007FF

// Word Address 0x00000258 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_ADR 32'h00000258
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_0_MSK 32'h0000003F

// Word Address 0x0000025C : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_ADR 32'h0000025C
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_1_MSK 32'h0000003F

// Word Address 0x00000260 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_ADR 32'h00000260
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_2_MSK 32'h0000003F

// Word Address 0x00000264 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_ADR 32'h00000264
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_3_MSK 32'h0000003F

// Word Address 0x00000268 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_ADR 32'h00000268
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_4_MSK 32'h0000003F

// Word Address 0x0000026C : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_ADR 32'h0000026C
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_5_MSK 32'h0000003F

// Word Address 0x00000270 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_ADR 32'h00000270
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_6_MSK 32'h0000003F

// Word Address 0x00000274 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_ADR 32'h00000274
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_7_MSK 32'h0000003F

// Word Address 0x00000278 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_ADR 32'h00000278
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_8_MSK 32'h0000003F

// Word Address 0x0000027C : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_ADR 32'h0000027C
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_9_MSK 32'h0000003F

// Word Address 0x00000280 : DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_ADR 32'h00000280
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M0_CFG_10_MSK 32'h0000003F

// Word Address 0x00000284 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_ADR 32'h00000284
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_0_MSK 32'h0000003F

// Word Address 0x00000288 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_ADR 32'h00000288
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_1_MSK 32'h0000003F

// Word Address 0x0000028C : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_ADR 32'h0000028C
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_2_MSK 32'h0000003F

// Word Address 0x00000290 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_ADR 32'h00000290
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_3_MSK 32'h0000003F

// Word Address 0x00000294 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_ADR 32'h00000294
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_4_MSK 32'h0000003F

// Word Address 0x00000298 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_ADR 32'h00000298
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_5_MSK 32'h0000003F

// Word Address 0x0000029C : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_ADR 32'h0000029C
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_6_MSK 32'h0000003F

// Word Address 0x000002A0 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_ADR 32'h000002A0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_7_MSK 32'h0000003F

// Word Address 0x000002A4 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_ADR 32'h000002A4
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_8_MSK 32'h0000003F

// Word Address 0x000002A8 : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_ADR 32'h000002A8
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_9_MSK 32'h0000003F

// Word Address 0x000002AC : DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10 (RW)
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_RANGE 5:0
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_WIDTH 6
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_ADR 32'h000002AC
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_POR 32'h00000001
`define DDR_CA_DQ_TX_EGRESS_ANA_M1_CFG_10_MSK 32'h0000003F

// Word Address 0x000002B0 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_ADR 32'h000002B0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_0_MSK 32'h0000007F

// Word Address 0x000002B4 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_ADR 32'h000002B4
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_1_MSK 32'h0000007F

// Word Address 0x000002B8 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_ADR 32'h000002B8
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_2_MSK 32'h0000007F

// Word Address 0x000002BC : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_ADR 32'h000002BC
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_3_MSK 32'h0000007F

// Word Address 0x000002C0 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_ADR 32'h000002C0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_4_MSK 32'h0000007F

// Word Address 0x000002C4 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_ADR 32'h000002C4
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_5_MSK 32'h0000007F

// Word Address 0x000002C8 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_ADR 32'h000002C8
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_6_MSK 32'h0000007F

// Word Address 0x000002CC : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_ADR 32'h000002CC
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_7_MSK 32'h0000007F

// Word Address 0x000002D0 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_ADR 32'h000002D0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_8_MSK 32'h0000007F

// Word Address 0x000002D4 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_ADR 32'h000002D4
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_9_MSK 32'h0000007F

// Word Address 0x000002D8 : DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_ADR 32'h000002D8
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M0_CFG_10_MSK 32'h0000007F

// Word Address 0x000002DC : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_ADR 32'h000002DC
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_0_MSK 32'h0000007F

// Word Address 0x000002E0 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_ADR 32'h000002E0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_1_MSK 32'h0000007F

// Word Address 0x000002E4 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_ADR 32'h000002E4
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_2_MSK 32'h0000007F

// Word Address 0x000002E8 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_ADR 32'h000002E8
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_3_MSK 32'h0000007F

// Word Address 0x000002EC : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_ADR 32'h000002EC
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_4_MSK 32'h0000007F

// Word Address 0x000002F0 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_ADR 32'h000002F0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_5_MSK 32'h0000007F

// Word Address 0x000002F4 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_ADR 32'h000002F4
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_6_MSK 32'h0000007F

// Word Address 0x000002F8 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_ADR 32'h000002F8
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_7_MSK 32'h0000007F

// Word Address 0x000002FC : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_ADR 32'h000002FC
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_8_MSK 32'h0000007F

// Word Address 0x00000300 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_ADR 32'h00000300
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_9_MSK 32'h0000007F

// Word Address 0x00000304 : DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10 (RW)
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_RANGE 6:0
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_WIDTH 7
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_ADR 32'h00000304
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_POR 32'h00000002
`define DDR_CA_DQ_TX_EGRESS_DIG_M1_CFG_10_MSK 32'h0000007F

// Word Address 0x00000308 : DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_ADR 32'h00000308
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_ODR_PI_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x0000030C : DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_ADR 32'h0000030C
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_ODR_PI_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000310 : DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_ADR 32'h00000310
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_ODR_PI_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000314 : DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_ADR 32'h00000314
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_ODR_PI_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000318 : DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_ADR 32'h00000318
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x0000031C : DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_ADR 32'h0000031C
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_0_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000320 : DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_ADR 32'h00000320
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000324 : DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_ADR 32'h00000324
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_0_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000328 : DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_ADR 32'h00000328
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x0000032C : DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_ADR 32'h0000032C
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_1_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000330 : DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_ADR 32'h00000330
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000334 : DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_ADR 32'h00000334
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_QDR_PI_1_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000338 : DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_ADR 32'h00000338
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x0000033C : DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_ADR 32'h0000033C
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_0_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000340 : DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_ADR 32'h00000340
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000344 : DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_ADR 32'h00000344
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_0_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000348 : DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_ADR 32'h00000348
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x0000034C : DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_ADR 32'h0000034C
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_1_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000350 : DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_ADR 32'h00000350
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000354 : DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_ADR 32'h00000354
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_DDR_PI_1_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000358 : DDR_CA_DQ_TX_PI_RT_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_ADR 32'h00000358
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_PI_RT_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x0000035C : DDR_CA_DQ_TX_PI_RT_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_ADR 32'h0000035C
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_PI_RT_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000360 : DDR_CA_DQ_TX_PI_RT_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_ADR 32'h00000360
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_PI_RT_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000364 : DDR_CA_DQ_TX_PI_RT_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_ADR 32'h00000364
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQ_TX_PI_RT_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000368 : DDR_CA_DQ_TX_RT_M0_R0_CFG (RW)
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_PIPE_EN_FIELD 10:0
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_PIPE_EN_FIELD_WIDTH 11
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_RANGE 10:0
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_WIDTH 11
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_ADR 32'h00000368
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_POR 32'h00000000
`define DDR_CA_DQ_TX_RT_M0_R0_CFG_MSK 32'h000007FF

// Word Address 0x0000036C : DDR_CA_DQ_TX_RT_M0_R1_CFG (RW)
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_PIPE_EN_FIELD 10:0
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_PIPE_EN_FIELD_WIDTH 11
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_RANGE 10:0
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_WIDTH 11
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_ADR 32'h0000036C
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_POR 32'h00000000
`define DDR_CA_DQ_TX_RT_M0_R1_CFG_MSK 32'h000007FF

// Word Address 0x00000370 : DDR_CA_DQ_TX_RT_M1_R0_CFG (RW)
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_PIPE_EN_FIELD 10:0
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_PIPE_EN_FIELD_WIDTH 11
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_RANGE 10:0
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_WIDTH 11
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_ADR 32'h00000370
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_POR 32'h00000000
`define DDR_CA_DQ_TX_RT_M1_R0_CFG_MSK 32'h000007FF

// Word Address 0x00000374 : DDR_CA_DQ_TX_RT_M1_R1_CFG (RW)
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_PIPE_EN_FIELD 10:0
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_PIPE_EN_FIELD_WIDTH 11
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_RANGE 10:0
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_WIDTH 11
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_ADR 32'h00000374
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_POR 32'h00000000
`define DDR_CA_DQ_TX_RT_M1_R1_CFG_MSK 32'h000007FF

// Word Address 0x00000378 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_ADR 32'h00000378
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_0_MSK 32'h000000FF

// Word Address 0x0000037C : DDR_CA_DQ_TX_SDR_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_ADR 32'h0000037C
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_1_MSK 32'h000000FF

// Word Address 0x00000380 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_ADR 32'h00000380
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_2_MSK 32'h000000FF

// Word Address 0x00000384 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_ADR 32'h00000384
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_3_MSK 32'h000000FF

// Word Address 0x00000388 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_ADR 32'h00000388
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_4_MSK 32'h000000FF

// Word Address 0x0000038C : DDR_CA_DQ_TX_SDR_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_ADR 32'h0000038C
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_5_MSK 32'h000000FF

// Word Address 0x00000390 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_ADR 32'h00000390
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_6_MSK 32'h000000FF

// Word Address 0x00000394 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_ADR 32'h00000394
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_7_MSK 32'h000000FF

// Word Address 0x00000398 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_ADR 32'h00000398
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_8_MSK 32'h000000FF

// Word Address 0x0000039C : DDR_CA_DQ_TX_SDR_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_ADR 32'h0000039C
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_9_MSK 32'h000000FF

// Word Address 0x000003A0 : DDR_CA_DQ_TX_SDR_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_ADR 32'h000003A0
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R0_CFG_10_MSK 32'h000000FF

// Word Address 0x000003A4 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_ADR 32'h000003A4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_0_MSK 32'h000000FF

// Word Address 0x000003A8 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_ADR 32'h000003A8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_1_MSK 32'h000000FF

// Word Address 0x000003AC : DDR_CA_DQ_TX_SDR_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_ADR 32'h000003AC
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_2_MSK 32'h000000FF

// Word Address 0x000003B0 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_ADR 32'h000003B0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_3_MSK 32'h000000FF

// Word Address 0x000003B4 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_ADR 32'h000003B4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_4_MSK 32'h000000FF

// Word Address 0x000003B8 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_ADR 32'h000003B8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_5_MSK 32'h000000FF

// Word Address 0x000003BC : DDR_CA_DQ_TX_SDR_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_ADR 32'h000003BC
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_6_MSK 32'h000000FF

// Word Address 0x000003C0 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_ADR 32'h000003C0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_7_MSK 32'h000000FF

// Word Address 0x000003C4 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_ADR 32'h000003C4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_8_MSK 32'h000000FF

// Word Address 0x000003C8 : DDR_CA_DQ_TX_SDR_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_ADR 32'h000003C8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_9_MSK 32'h000000FF

// Word Address 0x000003CC : DDR_CA_DQ_TX_SDR_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_ADR 32'h000003CC
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M0_R1_CFG_10_MSK 32'h000000FF

// Word Address 0x000003D0 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_ADR 32'h000003D0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_0_MSK 32'h000000FF

// Word Address 0x000003D4 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_ADR 32'h000003D4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_1_MSK 32'h000000FF

// Word Address 0x000003D8 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_ADR 32'h000003D8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_2_MSK 32'h000000FF

// Word Address 0x000003DC : DDR_CA_DQ_TX_SDR_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_ADR 32'h000003DC
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_3_MSK 32'h000000FF

// Word Address 0x000003E0 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_ADR 32'h000003E0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_4_MSK 32'h000000FF

// Word Address 0x000003E4 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_ADR 32'h000003E4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_5_MSK 32'h000000FF

// Word Address 0x000003E8 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_ADR 32'h000003E8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_6_MSK 32'h000000FF

// Word Address 0x000003EC : DDR_CA_DQ_TX_SDR_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_ADR 32'h000003EC
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_7_MSK 32'h000000FF

// Word Address 0x000003F0 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_ADR 32'h000003F0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_8_MSK 32'h000000FF

// Word Address 0x000003F4 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_ADR 32'h000003F4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_9_MSK 32'h000000FF

// Word Address 0x000003F8 : DDR_CA_DQ_TX_SDR_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_ADR 32'h000003F8
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R0_CFG_10_MSK 32'h000000FF

// Word Address 0x000003FC : DDR_CA_DQ_TX_SDR_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_ADR 32'h000003FC
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_0_MSK 32'h000000FF

// Word Address 0x00000400 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_ADR 32'h00000400
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_1_MSK 32'h000000FF

// Word Address 0x00000404 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_ADR 32'h00000404
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_2_MSK 32'h000000FF

// Word Address 0x00000408 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_ADR 32'h00000408
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_3_MSK 32'h000000FF

// Word Address 0x0000040C : DDR_CA_DQ_TX_SDR_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_ADR 32'h0000040C
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_4_MSK 32'h000000FF

// Word Address 0x00000410 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_ADR 32'h00000410
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_5_MSK 32'h000000FF

// Word Address 0x00000414 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_ADR 32'h00000414
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_6_MSK 32'h000000FF

// Word Address 0x00000418 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_ADR 32'h00000418
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_7_MSK 32'h000000FF

// Word Address 0x0000041C : DDR_CA_DQ_TX_SDR_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_ADR 32'h0000041C
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_8_MSK 32'h000000FF

// Word Address 0x00000420 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_ADR 32'h00000420
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_9_MSK 32'h000000FF

// Word Address 0x00000424 : DDR_CA_DQ_TX_SDR_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_RANGE 7:0
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_WIDTH 8
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_ADR 32'h00000424
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_M1_R1_CFG_10_MSK 32'h000000FF

// Word Address 0x00000428 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_ADR 32'h00000428
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_0_MSK 32'h77777777

// Word Address 0x0000042C : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_ADR 32'h0000042C
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_1_MSK 32'h77777777

// Word Address 0x00000430 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_ADR 32'h00000430
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_2_MSK 32'h77777777

// Word Address 0x00000434 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_ADR 32'h00000434
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_3_MSK 32'h77777777

// Word Address 0x00000438 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_ADR 32'h00000438
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_4_MSK 32'h77777777

// Word Address 0x0000043C : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_ADR 32'h0000043C
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_5_MSK 32'h77777777

// Word Address 0x00000440 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_ADR 32'h00000440
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_6_MSK 32'h77777777

// Word Address 0x00000444 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_ADR 32'h00000444
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_7_MSK 32'h77777777

// Word Address 0x00000448 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_ADR 32'h00000448
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_8_MSK 32'h77777777

// Word Address 0x0000044C : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_ADR 32'h0000044C
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_9_MSK 32'h77777777

// Word Address 0x00000450 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_ADR 32'h00000450
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R0_CFG_10_MSK 32'h77777777

// Word Address 0x00000454 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_ADR 32'h00000454
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_0_MSK 32'h77777777

// Word Address 0x00000458 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_ADR 32'h00000458
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_1_MSK 32'h77777777

// Word Address 0x0000045C : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_ADR 32'h0000045C
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_2_MSK 32'h77777777

// Word Address 0x00000460 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_ADR 32'h00000460
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_3_MSK 32'h77777777

// Word Address 0x00000464 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_ADR 32'h00000464
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_4_MSK 32'h77777777

// Word Address 0x00000468 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_ADR 32'h00000468
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_5_MSK 32'h77777777

// Word Address 0x0000046C : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_ADR 32'h0000046C
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_6_MSK 32'h77777777

// Word Address 0x00000470 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_ADR 32'h00000470
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_7_MSK 32'h77777777

// Word Address 0x00000474 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_ADR 32'h00000474
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_8_MSK 32'h77777777

// Word Address 0x00000478 : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_ADR 32'h00000478
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_9_MSK 32'h77777777

// Word Address 0x0000047C : DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_ADR 32'h0000047C
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M0_R1_CFG_10_MSK 32'h77777777

// Word Address 0x00000480 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_ADR 32'h00000480
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_0_MSK 32'h77777777

// Word Address 0x00000484 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_ADR 32'h00000484
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_1_MSK 32'h77777777

// Word Address 0x00000488 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_ADR 32'h00000488
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_2_MSK 32'h77777777

// Word Address 0x0000048C : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_ADR 32'h0000048C
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_3_MSK 32'h77777777

// Word Address 0x00000490 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_ADR 32'h00000490
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_4_MSK 32'h77777777

// Word Address 0x00000494 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_ADR 32'h00000494
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_5_MSK 32'h77777777

// Word Address 0x00000498 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_ADR 32'h00000498
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_6_MSK 32'h77777777

// Word Address 0x0000049C : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_ADR 32'h0000049C
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_7_MSK 32'h77777777

// Word Address 0x000004A0 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_ADR 32'h000004A0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_8_MSK 32'h77777777

// Word Address 0x000004A4 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_ADR 32'h000004A4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_9_MSK 32'h77777777

// Word Address 0x000004A8 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_ADR 32'h000004A8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R0_CFG_10_MSK 32'h77777777

// Word Address 0x000004AC : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_ADR 32'h000004AC
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_0_MSK 32'h77777777

// Word Address 0x000004B0 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_ADR 32'h000004B0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_1_MSK 32'h77777777

// Word Address 0x000004B4 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_ADR 32'h000004B4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_2_MSK 32'h77777777

// Word Address 0x000004B8 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_ADR 32'h000004B8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_3_MSK 32'h77777777

// Word Address 0x000004BC : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_ADR 32'h000004BC
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_4_MSK 32'h77777777

// Word Address 0x000004C0 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_ADR 32'h000004C0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_5_MSK 32'h77777777

// Word Address 0x000004C4 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_ADR 32'h000004C4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_6_MSK 32'h77777777

// Word Address 0x000004C8 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_ADR 32'h000004C8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_7_MSK 32'h77777777

// Word Address 0x000004CC : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_ADR 32'h000004CC
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_8_MSK 32'h77777777

// Word Address 0x000004D0 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_ADR 32'h000004D0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_9_MSK 32'h77777777

// Word Address 0x000004D4 : DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_RANGE 30:0
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_WIDTH 31
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_ADR 32'h000004D4
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_X_SEL_M1_R1_CFG_10_MSK 32'h77777777

// Word Address 0x000004D8 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_ADR 32'h000004D8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0_MSK 32'h33333333

// Word Address 0x000004DC : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_ADR 32'h000004DC
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1_MSK 32'h33333333

// Word Address 0x000004E0 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_ADR 32'h000004E0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2_MSK 32'h33333333

// Word Address 0x000004E4 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_ADR 32'h000004E4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3_MSK 32'h33333333

// Word Address 0x000004E8 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_ADR 32'h000004E8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4_MSK 32'h33333333

// Word Address 0x000004EC : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_ADR 32'h000004EC
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5_MSK 32'h33333333

// Word Address 0x000004F0 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_ADR 32'h000004F0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6_MSK 32'h33333333

// Word Address 0x000004F4 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_ADR 32'h000004F4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7_MSK 32'h33333333

// Word Address 0x000004F8 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_ADR 32'h000004F8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8_MSK 32'h33333333

// Word Address 0x000004FC : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_ADR 32'h000004FC
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9_MSK 32'h33333333

// Word Address 0x00000500 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_ADR 32'h00000500
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10_MSK 32'h33333333

// Word Address 0x00000504 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_ADR 32'h00000504
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0_MSK 32'h33333333

// Word Address 0x00000508 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_ADR 32'h00000508
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1_MSK 32'h33333333

// Word Address 0x0000050C : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_ADR 32'h0000050C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2_MSK 32'h33333333

// Word Address 0x00000510 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_ADR 32'h00000510
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3_MSK 32'h33333333

// Word Address 0x00000514 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_ADR 32'h00000514
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4_MSK 32'h33333333

// Word Address 0x00000518 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_ADR 32'h00000518
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5_MSK 32'h33333333

// Word Address 0x0000051C : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_ADR 32'h0000051C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6_MSK 32'h33333333

// Word Address 0x00000520 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_ADR 32'h00000520
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7_MSK 32'h33333333

// Word Address 0x00000524 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_ADR 32'h00000524
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8_MSK 32'h33333333

// Word Address 0x00000528 : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_ADR 32'h00000528
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9_MSK 32'h33333333

// Word Address 0x0000052C : DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_ADR 32'h0000052C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10_MSK 32'h33333333

// Word Address 0x00000530 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_ADR 32'h00000530
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0_MSK 32'h33333333

// Word Address 0x00000534 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_ADR 32'h00000534
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1_MSK 32'h33333333

// Word Address 0x00000538 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_ADR 32'h00000538
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2_MSK 32'h33333333

// Word Address 0x0000053C : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_ADR 32'h0000053C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3_MSK 32'h33333333

// Word Address 0x00000540 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_ADR 32'h00000540
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4_MSK 32'h33333333

// Word Address 0x00000544 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_ADR 32'h00000544
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5_MSK 32'h33333333

// Word Address 0x00000548 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_ADR 32'h00000548
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6_MSK 32'h33333333

// Word Address 0x0000054C : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_ADR 32'h0000054C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7_MSK 32'h33333333

// Word Address 0x00000550 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_ADR 32'h00000550
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8_MSK 32'h33333333

// Word Address 0x00000554 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_ADR 32'h00000554
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9_MSK 32'h33333333

// Word Address 0x00000558 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_ADR 32'h00000558
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10_MSK 32'h33333333

// Word Address 0x0000055C : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_ADR 32'h0000055C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0_MSK 32'h33333333

// Word Address 0x00000560 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_ADR 32'h00000560
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1_MSK 32'h33333333

// Word Address 0x00000564 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_ADR 32'h00000564
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2_MSK 32'h33333333

// Word Address 0x00000568 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_ADR 32'h00000568
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3_MSK 32'h33333333

// Word Address 0x0000056C : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_ADR 32'h0000056C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4_MSK 32'h33333333

// Word Address 0x00000570 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_ADR 32'h00000570
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5_MSK 32'h33333333

// Word Address 0x00000574 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_ADR 32'h00000574
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6_MSK 32'h33333333

// Word Address 0x00000578 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_ADR 32'h00000578
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7_MSK 32'h33333333

// Word Address 0x0000057C : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_ADR 32'h0000057C
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8_MSK 32'h33333333

// Word Address 0x00000580 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_ADR 32'h00000580
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9_MSK 32'h33333333

// Word Address 0x00000584 : DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P0_FIELD 1:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P1_FIELD 5:4
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P2_FIELD 9:8
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P3_FIELD 13:12
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P4_FIELD 17:16
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P5_FIELD 21:20
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P6_FIELD 25:24
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P7_FIELD 29:28
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_RANGE 29:0
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_WIDTH 30
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_ADR 32'h00000584
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10_MSK 32'h33333333

// Word Address 0x00000588 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_ADR 32'h00000588
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_0_MSK 32'h0000000F

// Word Address 0x0000058C : DDR_CA_DQ_TX_DDR_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_ADR 32'h0000058C
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_1_MSK 32'h0000000F

// Word Address 0x00000590 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_ADR 32'h00000590
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_2_MSK 32'h0000000F

// Word Address 0x00000594 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_ADR 32'h00000594
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_3_MSK 32'h0000000F

// Word Address 0x00000598 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_ADR 32'h00000598
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_4_MSK 32'h0000000F

// Word Address 0x0000059C : DDR_CA_DQ_TX_DDR_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_ADR 32'h0000059C
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_5_MSK 32'h0000000F

// Word Address 0x000005A0 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_ADR 32'h000005A0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_6_MSK 32'h0000000F

// Word Address 0x000005A4 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_ADR 32'h000005A4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_7_MSK 32'h0000000F

// Word Address 0x000005A8 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_ADR 32'h000005A8
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_8_MSK 32'h0000000F

// Word Address 0x000005AC : DDR_CA_DQ_TX_DDR_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_ADR 32'h000005AC
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_9_MSK 32'h0000000F

// Word Address 0x000005B0 : DDR_CA_DQ_TX_DDR_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_ADR 32'h000005B0
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R0_CFG_10_MSK 32'h0000000F

// Word Address 0x000005B4 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_ADR 32'h000005B4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_0_MSK 32'h0000000F

// Word Address 0x000005B8 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_ADR 32'h000005B8
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_1_MSK 32'h0000000F

// Word Address 0x000005BC : DDR_CA_DQ_TX_DDR_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_ADR 32'h000005BC
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_2_MSK 32'h0000000F

// Word Address 0x000005C0 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_ADR 32'h000005C0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_3_MSK 32'h0000000F

// Word Address 0x000005C4 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_ADR 32'h000005C4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_4_MSK 32'h0000000F

// Word Address 0x000005C8 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_ADR 32'h000005C8
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_5_MSK 32'h0000000F

// Word Address 0x000005CC : DDR_CA_DQ_TX_DDR_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_ADR 32'h000005CC
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_6_MSK 32'h0000000F

// Word Address 0x000005D0 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_ADR 32'h000005D0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_7_MSK 32'h0000000F

// Word Address 0x000005D4 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_ADR 32'h000005D4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_8_MSK 32'h0000000F

// Word Address 0x000005D8 : DDR_CA_DQ_TX_DDR_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_ADR 32'h000005D8
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_9_MSK 32'h0000000F

// Word Address 0x000005DC : DDR_CA_DQ_TX_DDR_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_ADR 32'h000005DC
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M0_R1_CFG_10_MSK 32'h0000000F

// Word Address 0x000005E0 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_ADR 32'h000005E0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_0_MSK 32'h0000000F

// Word Address 0x000005E4 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_ADR 32'h000005E4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_1_MSK 32'h0000000F

// Word Address 0x000005E8 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_ADR 32'h000005E8
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_2_MSK 32'h0000000F

// Word Address 0x000005EC : DDR_CA_DQ_TX_DDR_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_ADR 32'h000005EC
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_3_MSK 32'h0000000F

// Word Address 0x000005F0 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_ADR 32'h000005F0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_4_MSK 32'h0000000F

// Word Address 0x000005F4 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_ADR 32'h000005F4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_5_MSK 32'h0000000F

// Word Address 0x000005F8 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_ADR 32'h000005F8
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_6_MSK 32'h0000000F

// Word Address 0x000005FC : DDR_CA_DQ_TX_DDR_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_ADR 32'h000005FC
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_7_MSK 32'h0000000F

// Word Address 0x00000600 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_ADR 32'h00000600
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_8_MSK 32'h0000000F

// Word Address 0x00000604 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_ADR 32'h00000604
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_9_MSK 32'h0000000F

// Word Address 0x00000608 : DDR_CA_DQ_TX_DDR_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_ADR 32'h00000608
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R0_CFG_10_MSK 32'h0000000F

// Word Address 0x0000060C : DDR_CA_DQ_TX_DDR_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_ADR 32'h0000060C
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_0_MSK 32'h0000000F

// Word Address 0x00000610 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_ADR 32'h00000610
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_1_MSK 32'h0000000F

// Word Address 0x00000614 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_ADR 32'h00000614
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_2_MSK 32'h0000000F

// Word Address 0x00000618 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_ADR 32'h00000618
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_3_MSK 32'h0000000F

// Word Address 0x0000061C : DDR_CA_DQ_TX_DDR_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_ADR 32'h0000061C
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_4_MSK 32'h0000000F

// Word Address 0x00000620 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_ADR 32'h00000620
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_5_MSK 32'h0000000F

// Word Address 0x00000624 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_ADR 32'h00000624
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_6_MSK 32'h0000000F

// Word Address 0x00000628 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_ADR 32'h00000628
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_7_MSK 32'h0000000F

// Word Address 0x0000062C : DDR_CA_DQ_TX_DDR_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_ADR 32'h0000062C
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_8_MSK 32'h0000000F

// Word Address 0x00000630 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_ADR 32'h00000630
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_9_MSK 32'h0000000F

// Word Address 0x00000634 : DDR_CA_DQ_TX_DDR_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_RANGE 3:0
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_WIDTH 4
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_ADR 32'h00000634
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_M1_R1_CFG_10_MSK 32'h0000000F

// Word Address 0x00000638 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_ADR 32'h00000638
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_0_MSK 32'h00003333

// Word Address 0x0000063C : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_ADR 32'h0000063C
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_1_MSK 32'h00003333

// Word Address 0x00000640 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_ADR 32'h00000640
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_2_MSK 32'h00003333

// Word Address 0x00000644 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_ADR 32'h00000644
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_3_MSK 32'h00003333

// Word Address 0x00000648 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_ADR 32'h00000648
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_4_MSK 32'h00003333

// Word Address 0x0000064C : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_ADR 32'h0000064C
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_5_MSK 32'h00003333

// Word Address 0x00000650 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_ADR 32'h00000650
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_6_MSK 32'h00003333

// Word Address 0x00000654 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_ADR 32'h00000654
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_7_MSK 32'h00003333

// Word Address 0x00000658 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_ADR 32'h00000658
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_8_MSK 32'h00003333

// Word Address 0x0000065C : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_ADR 32'h0000065C
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_9_MSK 32'h00003333

// Word Address 0x00000660 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_ADR 32'h00000660
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R0_CFG_10_MSK 32'h00003333

// Word Address 0x00000664 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_ADR 32'h00000664
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_0_MSK 32'h00003333

// Word Address 0x00000668 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_ADR 32'h00000668
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_1_MSK 32'h00003333

// Word Address 0x0000066C : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_ADR 32'h0000066C
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_2_MSK 32'h00003333

// Word Address 0x00000670 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_ADR 32'h00000670
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_3_MSK 32'h00003333

// Word Address 0x00000674 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_ADR 32'h00000674
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_4_MSK 32'h00003333

// Word Address 0x00000678 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_ADR 32'h00000678
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_5_MSK 32'h00003333

// Word Address 0x0000067C : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_ADR 32'h0000067C
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_6_MSK 32'h00003333

// Word Address 0x00000680 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_ADR 32'h00000680
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_7_MSK 32'h00003333

// Word Address 0x00000684 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_ADR 32'h00000684
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_8_MSK 32'h00003333

// Word Address 0x00000688 : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_ADR 32'h00000688
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_9_MSK 32'h00003333

// Word Address 0x0000068C : DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_ADR 32'h0000068C
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M0_R1_CFG_10_MSK 32'h00003333

// Word Address 0x00000690 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_ADR 32'h00000690
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_0_MSK 32'h00003333

// Word Address 0x00000694 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_ADR 32'h00000694
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_1_MSK 32'h00003333

// Word Address 0x00000698 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_ADR 32'h00000698
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_2_MSK 32'h00003333

// Word Address 0x0000069C : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_ADR 32'h0000069C
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_3_MSK 32'h00003333

// Word Address 0x000006A0 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_ADR 32'h000006A0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_4_MSK 32'h00003333

// Word Address 0x000006A4 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_ADR 32'h000006A4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_5_MSK 32'h00003333

// Word Address 0x000006A8 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_ADR 32'h000006A8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_6_MSK 32'h00003333

// Word Address 0x000006AC : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_ADR 32'h000006AC
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_7_MSK 32'h00003333

// Word Address 0x000006B0 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_ADR 32'h000006B0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_8_MSK 32'h00003333

// Word Address 0x000006B4 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_ADR 32'h000006B4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_9_MSK 32'h00003333

// Word Address 0x000006B8 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_ADR 32'h000006B8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R0_CFG_10_MSK 32'h00003333

// Word Address 0x000006BC : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_ADR 32'h000006BC
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_0_MSK 32'h00003333

// Word Address 0x000006C0 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_ADR 32'h000006C0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_1_MSK 32'h00003333

// Word Address 0x000006C4 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_ADR 32'h000006C4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_2_MSK 32'h00003333

// Word Address 0x000006C8 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_ADR 32'h000006C8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_3_MSK 32'h00003333

// Word Address 0x000006CC : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_ADR 32'h000006CC
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_4_MSK 32'h00003333

// Word Address 0x000006D0 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_ADR 32'h000006D0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_5_MSK 32'h00003333

// Word Address 0x000006D4 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_ADR 32'h000006D4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_6_MSK 32'h00003333

// Word Address 0x000006D8 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_ADR 32'h000006D8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_7_MSK 32'h00003333

// Word Address 0x000006DC : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_ADR 32'h000006DC
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_8_MSK 32'h00003333

// Word Address 0x000006E0 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_ADR 32'h000006E0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_9_MSK 32'h00003333

// Word Address 0x000006E4 : DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_RANGE 13:0
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_WIDTH 14
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_ADR 32'h000006E4
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_DDR_X_SEL_M1_R1_CFG_10_MSK 32'h00003333

// Word Address 0x000006E8 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_ADR 32'h000006E8
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_0_MSK 32'h00000003

// Word Address 0x000006EC : DDR_CA_DQ_TX_QDR_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_ADR 32'h000006EC
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_1_MSK 32'h00000003

// Word Address 0x000006F0 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_ADR 32'h000006F0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_2_MSK 32'h00000003

// Word Address 0x000006F4 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_ADR 32'h000006F4
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_3_MSK 32'h00000003

// Word Address 0x000006F8 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_ADR 32'h000006F8
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_4_MSK 32'h00000003

// Word Address 0x000006FC : DDR_CA_DQ_TX_QDR_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_ADR 32'h000006FC
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_5_MSK 32'h00000003

// Word Address 0x00000700 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_ADR 32'h00000700
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_6_MSK 32'h00000003

// Word Address 0x00000704 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_ADR 32'h00000704
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_7_MSK 32'h00000003

// Word Address 0x00000708 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_ADR 32'h00000708
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_8_MSK 32'h00000003

// Word Address 0x0000070C : DDR_CA_DQ_TX_QDR_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_ADR 32'h0000070C
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_9_MSK 32'h00000003

// Word Address 0x00000710 : DDR_CA_DQ_TX_QDR_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_ADR 32'h00000710
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R0_CFG_10_MSK 32'h00000003

// Word Address 0x00000714 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_ADR 32'h00000714
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_0_MSK 32'h00000003

// Word Address 0x00000718 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_ADR 32'h00000718
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_1_MSK 32'h00000003

// Word Address 0x0000071C : DDR_CA_DQ_TX_QDR_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_ADR 32'h0000071C
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_2_MSK 32'h00000003

// Word Address 0x00000720 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_ADR 32'h00000720
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_3_MSK 32'h00000003

// Word Address 0x00000724 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_ADR 32'h00000724
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_4_MSK 32'h00000003

// Word Address 0x00000728 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_ADR 32'h00000728
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_5_MSK 32'h00000003

// Word Address 0x0000072C : DDR_CA_DQ_TX_QDR_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_ADR 32'h0000072C
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_6_MSK 32'h00000003

// Word Address 0x00000730 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_ADR 32'h00000730
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_7_MSK 32'h00000003

// Word Address 0x00000734 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_ADR 32'h00000734
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_8_MSK 32'h00000003

// Word Address 0x00000738 : DDR_CA_DQ_TX_QDR_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_ADR 32'h00000738
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_9_MSK 32'h00000003

// Word Address 0x0000073C : DDR_CA_DQ_TX_QDR_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_ADR 32'h0000073C
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M0_R1_CFG_10_MSK 32'h00000003

// Word Address 0x00000740 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_ADR 32'h00000740
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_0_MSK 32'h00000003

// Word Address 0x00000744 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_ADR 32'h00000744
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_1_MSK 32'h00000003

// Word Address 0x00000748 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_ADR 32'h00000748
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_2_MSK 32'h00000003

// Word Address 0x0000074C : DDR_CA_DQ_TX_QDR_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_ADR 32'h0000074C
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_3_MSK 32'h00000003

// Word Address 0x00000750 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_ADR 32'h00000750
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_4_MSK 32'h00000003

// Word Address 0x00000754 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_ADR 32'h00000754
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_5_MSK 32'h00000003

// Word Address 0x00000758 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_ADR 32'h00000758
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_6_MSK 32'h00000003

// Word Address 0x0000075C : DDR_CA_DQ_TX_QDR_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_ADR 32'h0000075C
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_7_MSK 32'h00000003

// Word Address 0x00000760 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_ADR 32'h00000760
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_8_MSK 32'h00000003

// Word Address 0x00000764 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_ADR 32'h00000764
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_9_MSK 32'h00000003

// Word Address 0x00000768 : DDR_CA_DQ_TX_QDR_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_ADR 32'h00000768
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R0_CFG_10_MSK 32'h00000003

// Word Address 0x0000076C : DDR_CA_DQ_TX_QDR_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_ADR 32'h0000076C
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_0_MSK 32'h00000003

// Word Address 0x00000770 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_ADR 32'h00000770
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_1_MSK 32'h00000003

// Word Address 0x00000774 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_ADR 32'h00000774
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_2_MSK 32'h00000003

// Word Address 0x00000778 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_ADR 32'h00000778
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_3_MSK 32'h00000003

// Word Address 0x0000077C : DDR_CA_DQ_TX_QDR_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_ADR 32'h0000077C
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_4_MSK 32'h00000003

// Word Address 0x00000780 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_ADR 32'h00000780
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_5_MSK 32'h00000003

// Word Address 0x00000784 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_ADR 32'h00000784
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_6_MSK 32'h00000003

// Word Address 0x00000788 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_ADR 32'h00000788
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_7_MSK 32'h00000003

// Word Address 0x0000078C : DDR_CA_DQ_TX_QDR_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_ADR 32'h0000078C
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_8_MSK 32'h00000003

// Word Address 0x00000790 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_ADR 32'h00000790
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_9_MSK 32'h00000003

// Word Address 0x00000794 : DDR_CA_DQ_TX_QDR_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_RANGE 1:0
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_WIDTH 2
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_ADR 32'h00000794
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_M1_R1_CFG_10_MSK 32'h00000003

// Word Address 0x00000798 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_ADR 32'h00000798
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_0_MSK 32'h00000011

// Word Address 0x0000079C : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_ADR 32'h0000079C
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_1_MSK 32'h00000011

// Word Address 0x000007A0 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_ADR 32'h000007A0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_2_MSK 32'h00000011

// Word Address 0x000007A4 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_ADR 32'h000007A4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_3_MSK 32'h00000011

// Word Address 0x000007A8 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_ADR 32'h000007A8
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_4_MSK 32'h00000011

// Word Address 0x000007AC : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_ADR 32'h000007AC
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_5_MSK 32'h00000011

// Word Address 0x000007B0 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_ADR 32'h000007B0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_6_MSK 32'h00000011

// Word Address 0x000007B4 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_ADR 32'h000007B4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_7_MSK 32'h00000011

// Word Address 0x000007B8 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_ADR 32'h000007B8
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_8_MSK 32'h00000011

// Word Address 0x000007BC : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_ADR 32'h000007BC
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_9_MSK 32'h00000011

// Word Address 0x000007C0 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_ADR 32'h000007C0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R0_CFG_10_MSK 32'h00000011

// Word Address 0x000007C4 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_ADR 32'h000007C4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_0_MSK 32'h00000011

// Word Address 0x000007C8 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_ADR 32'h000007C8
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_1_MSK 32'h00000011

// Word Address 0x000007CC : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_ADR 32'h000007CC
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_2_MSK 32'h00000011

// Word Address 0x000007D0 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_ADR 32'h000007D0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_3_MSK 32'h00000011

// Word Address 0x000007D4 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_ADR 32'h000007D4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_4_MSK 32'h00000011

// Word Address 0x000007D8 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_ADR 32'h000007D8
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_5_MSK 32'h00000011

// Word Address 0x000007DC : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_ADR 32'h000007DC
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_6_MSK 32'h00000011

// Word Address 0x000007E0 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_ADR 32'h000007E0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_7_MSK 32'h00000011

// Word Address 0x000007E4 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_ADR 32'h000007E4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_8_MSK 32'h00000011

// Word Address 0x000007E8 : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_ADR 32'h000007E8
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_9_MSK 32'h00000011

// Word Address 0x000007EC : DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_ADR 32'h000007EC
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M0_R1_CFG_10_MSK 32'h00000011

// Word Address 0x000007F0 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_ADR 32'h000007F0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_0_MSK 32'h00000011

// Word Address 0x000007F4 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_ADR 32'h000007F4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_1_MSK 32'h00000011

// Word Address 0x000007F8 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_ADR 32'h000007F8
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_2_MSK 32'h00000011

// Word Address 0x000007FC : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_ADR 32'h000007FC
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_3_MSK 32'h00000011

// Word Address 0x00000800 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_ADR 32'h00000800
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_4_MSK 32'h00000011

// Word Address 0x00000804 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_ADR 32'h00000804
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_5_MSK 32'h00000011

// Word Address 0x00000808 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_ADR 32'h00000808
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_6_MSK 32'h00000011

// Word Address 0x0000080C : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_ADR 32'h0000080C
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_7_MSK 32'h00000011

// Word Address 0x00000810 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_ADR 32'h00000810
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_8_MSK 32'h00000011

// Word Address 0x00000814 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_ADR 32'h00000814
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_9_MSK 32'h00000011

// Word Address 0x00000818 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_ADR 32'h00000818
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R0_CFG_10_MSK 32'h00000011

// Word Address 0x0000081C : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_ADR 32'h0000081C
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_0_MSK 32'h00000011

// Word Address 0x00000820 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_ADR 32'h00000820
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_1_MSK 32'h00000011

// Word Address 0x00000824 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_ADR 32'h00000824
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_2_MSK 32'h00000011

// Word Address 0x00000828 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_ADR 32'h00000828
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_3_MSK 32'h00000011

// Word Address 0x0000082C : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_ADR 32'h0000082C
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_4_MSK 32'h00000011

// Word Address 0x00000830 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_ADR 32'h00000830
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_5_MSK 32'h00000011

// Word Address 0x00000834 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_ADR 32'h00000834
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_6_MSK 32'h00000011

// Word Address 0x00000838 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_ADR 32'h00000838
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_7_MSK 32'h00000011

// Word Address 0x0000083C : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_ADR 32'h0000083C
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_8_MSK 32'h00000011

// Word Address 0x00000840 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_ADR 32'h00000840
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_9_MSK 32'h00000011

// Word Address 0x00000844 : DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_X_SEL_P0_FIELD 0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_X_SEL_P1_FIELD 4
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_RANGE 4:0
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_WIDTH 5
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_ADR 32'h00000844
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_POR 32'h00000000
`define DDR_CA_DQ_TX_QDR_X_SEL_M1_R1_CFG_10_MSK 32'h00000011

// Word Address 0x00000848 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_ADR 32'h00000848
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_0_MSK 32'h000001FF

// Word Address 0x0000084C : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_ADR 32'h0000084C
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_1_MSK 32'h000001FF

// Word Address 0x00000850 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_ADR 32'h00000850
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_2_MSK 32'h000001FF

// Word Address 0x00000854 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_ADR 32'h00000854
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_3_MSK 32'h000001FF

// Word Address 0x00000858 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_ADR 32'h00000858
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_4_MSK 32'h000001FF

// Word Address 0x0000085C : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_ADR 32'h0000085C
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_5_MSK 32'h000001FF

// Word Address 0x00000860 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_ADR 32'h00000860
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_6_MSK 32'h000001FF

// Word Address 0x00000864 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_ADR 32'h00000864
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_7_MSK 32'h000001FF

// Word Address 0x00000868 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_ADR 32'h00000868
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_8_MSK 32'h000001FF

// Word Address 0x0000086C : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_ADR 32'h0000086C
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_9_MSK 32'h000001FF

// Word Address 0x00000870 : DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_ADR 32'h00000870
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R0_CFG_10_MSK 32'h000001FF

// Word Address 0x00000874 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_ADR 32'h00000874
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_0_MSK 32'h000001FF

// Word Address 0x00000878 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_ADR 32'h00000878
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_1_MSK 32'h000001FF

// Word Address 0x0000087C : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_ADR 32'h0000087C
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_2_MSK 32'h000001FF

// Word Address 0x00000880 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_ADR 32'h00000880
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_3_MSK 32'h000001FF

// Word Address 0x00000884 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_ADR 32'h00000884
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_4_MSK 32'h000001FF

// Word Address 0x00000888 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_ADR 32'h00000888
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_5_MSK 32'h000001FF

// Word Address 0x0000088C : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_ADR 32'h0000088C
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_6_MSK 32'h000001FF

// Word Address 0x00000890 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_ADR 32'h00000890
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_7_MSK 32'h000001FF

// Word Address 0x00000894 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_ADR 32'h00000894
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_8_MSK 32'h000001FF

// Word Address 0x00000898 : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_ADR 32'h00000898
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_9_MSK 32'h000001FF

// Word Address 0x0000089C : DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_ADR 32'h0000089C
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M0_R1_CFG_10_MSK 32'h000001FF

// Word Address 0x000008A0 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_ADR 32'h000008A0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_0_MSK 32'h000001FF

// Word Address 0x000008A4 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_ADR 32'h000008A4
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_1_MSK 32'h000001FF

// Word Address 0x000008A8 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_ADR 32'h000008A8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_2_MSK 32'h000001FF

// Word Address 0x000008AC : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_ADR 32'h000008AC
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_3_MSK 32'h000001FF

// Word Address 0x000008B0 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_ADR 32'h000008B0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_4_MSK 32'h000001FF

// Word Address 0x000008B4 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_ADR 32'h000008B4
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_5_MSK 32'h000001FF

// Word Address 0x000008B8 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_ADR 32'h000008B8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_6_MSK 32'h000001FF

// Word Address 0x000008BC : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_ADR 32'h000008BC
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_7_MSK 32'h000001FF

// Word Address 0x000008C0 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_ADR 32'h000008C0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_8_MSK 32'h000001FF

// Word Address 0x000008C4 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_ADR 32'h000008C4
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_9_MSK 32'h000001FF

// Word Address 0x000008C8 : DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_ADR 32'h000008C8
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R0_CFG_10_MSK 32'h000001FF

// Word Address 0x000008CC : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_ADR 32'h000008CC
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_0_MSK 32'h000001FF

// Word Address 0x000008D0 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_ADR 32'h000008D0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_1_MSK 32'h000001FF

// Word Address 0x000008D4 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_ADR 32'h000008D4
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_2_MSK 32'h000001FF

// Word Address 0x000008D8 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_ADR 32'h000008D8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_3_MSK 32'h000001FF

// Word Address 0x000008DC : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_ADR 32'h000008DC
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_4_MSK 32'h000001FF

// Word Address 0x000008E0 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_ADR 32'h000008E0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_5_MSK 32'h000001FF

// Word Address 0x000008E4 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_ADR 32'h000008E4
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_6_MSK 32'h000001FF

// Word Address 0x000008E8 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_ADR 32'h000008E8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_7_MSK 32'h000001FF

// Word Address 0x000008EC : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_ADR 32'h000008EC
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_8_MSK 32'h000001FF

// Word Address 0x000008F0 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_ADR 32'h000008F0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_9_MSK 32'h000001FF

// Word Address 0x000008F4 : DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10 (RW)
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_EN_FIELD 8
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_EN_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_GEAR_FIELD 7:6
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_RANGE 8:0
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_WIDTH 9
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_ADR 32'h000008F4
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_POR 32'h00000100
`define DDR_CA_DQ_TX_LPDE_M1_R1_CFG_10_MSK 32'h000001FF

// Word Address 0x000008F8 : DDR_CA_DQ_TX_IO_M0_CFG_0 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_0_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_0_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_0_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_0_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_0_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_0_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_0_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_0_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_0_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_0_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_0_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_0_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_0_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_0_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_0_ADR 32'h000008F8
`define DDR_CA_DQ_TX_IO_M0_CFG_0_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_0_MSK 32'h00000FFF

// Word Address 0x000008FC : DDR_CA_DQ_TX_IO_M0_CFG_1 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_1_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_1_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_1_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_1_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_1_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_1_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_1_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_1_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_1_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_1_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_1_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_1_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_1_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_1_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_1_ADR 32'h000008FC
`define DDR_CA_DQ_TX_IO_M0_CFG_1_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_1_MSK 32'h00000FFF

// Word Address 0x00000900 : DDR_CA_DQ_TX_IO_M0_CFG_2 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_2_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_2_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_2_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_2_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_2_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_2_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_2_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_2_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_2_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_2_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_2_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_2_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_2_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_2_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_2_ADR 32'h00000900
`define DDR_CA_DQ_TX_IO_M0_CFG_2_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_2_MSK 32'h00000FFF

// Word Address 0x00000904 : DDR_CA_DQ_TX_IO_M0_CFG_3 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_3_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_3_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_3_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_3_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_3_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_3_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_3_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_3_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_3_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_3_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_3_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_3_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_3_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_3_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_3_ADR 32'h00000904
`define DDR_CA_DQ_TX_IO_M0_CFG_3_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_3_MSK 32'h00000FFF

// Word Address 0x00000908 : DDR_CA_DQ_TX_IO_M0_CFG_4 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_4_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_4_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_4_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_4_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_4_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_4_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_4_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_4_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_4_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_4_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_4_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_4_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_4_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_4_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_4_ADR 32'h00000908
`define DDR_CA_DQ_TX_IO_M0_CFG_4_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_4_MSK 32'h00000FFF

// Word Address 0x0000090C : DDR_CA_DQ_TX_IO_M0_CFG_5 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_5_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_5_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_5_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_5_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_5_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_5_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_5_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_5_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_5_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_5_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_5_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_5_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_5_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_5_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_5_ADR 32'h0000090C
`define DDR_CA_DQ_TX_IO_M0_CFG_5_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_5_MSK 32'h00000FFF

// Word Address 0x00000910 : DDR_CA_DQ_TX_IO_M0_CFG_6 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_6_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_6_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_6_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_6_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_6_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_6_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_6_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_6_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_6_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_6_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_6_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_6_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_6_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_6_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_6_ADR 32'h00000910
`define DDR_CA_DQ_TX_IO_M0_CFG_6_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_6_MSK 32'h00000FFF

// Word Address 0x00000914 : DDR_CA_DQ_TX_IO_M0_CFG_7 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_7_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_7_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_7_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_7_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_7_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_7_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_7_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_7_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_7_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_7_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_7_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_7_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_7_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_7_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_7_ADR 32'h00000914
`define DDR_CA_DQ_TX_IO_M0_CFG_7_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_7_MSK 32'h00000FFF

// Word Address 0x00000918 : DDR_CA_DQ_TX_IO_M0_CFG_8 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_8_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_8_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_8_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_8_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_8_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_8_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_8_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_8_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_8_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_8_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_8_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_8_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_8_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_8_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_8_ADR 32'h00000918
`define DDR_CA_DQ_TX_IO_M0_CFG_8_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_8_MSK 32'h00000FFF

// Word Address 0x0000091C : DDR_CA_DQ_TX_IO_M0_CFG_9 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_9_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_9_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_9_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_9_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_9_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_9_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_9_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_9_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_9_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_9_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_9_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_9_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_9_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_9_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_9_ADR 32'h0000091C
`define DDR_CA_DQ_TX_IO_M0_CFG_9_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_9_MSK 32'h00000FFF

// Word Address 0x00000920 : DDR_CA_DQ_TX_IO_M0_CFG_10 (RW)
`define DDR_CA_DQ_TX_IO_M0_CFG_10_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M0_CFG_10_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_10_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M0_CFG_10_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_10_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M0_CFG_10_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_10_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M0_CFG_10_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_10_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M0_CFG_10_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M0_CFG_10_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M0_CFG_10_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M0_CFG_10_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M0_CFG_10_WIDTH 12
`define DDR_CA_DQ_TX_IO_M0_CFG_10_ADR 32'h00000920
`define DDR_CA_DQ_TX_IO_M0_CFG_10_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M0_CFG_10_MSK 32'h00000FFF

// Word Address 0x00000924 : DDR_CA_DQ_TX_IO_M1_CFG_0 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_0_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_0_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_0_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_0_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_0_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_0_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_0_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_0_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_0_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_0_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_0_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_0_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_0_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_0_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_0_ADR 32'h00000924
`define DDR_CA_DQ_TX_IO_M1_CFG_0_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_0_MSK 32'h00000FFF

// Word Address 0x00000928 : DDR_CA_DQ_TX_IO_M1_CFG_1 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_1_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_1_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_1_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_1_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_1_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_1_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_1_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_1_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_1_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_1_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_1_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_1_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_1_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_1_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_1_ADR 32'h00000928
`define DDR_CA_DQ_TX_IO_M1_CFG_1_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_1_MSK 32'h00000FFF

// Word Address 0x0000092C : DDR_CA_DQ_TX_IO_M1_CFG_2 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_2_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_2_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_2_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_2_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_2_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_2_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_2_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_2_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_2_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_2_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_2_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_2_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_2_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_2_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_2_ADR 32'h0000092C
`define DDR_CA_DQ_TX_IO_M1_CFG_2_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_2_MSK 32'h00000FFF

// Word Address 0x00000930 : DDR_CA_DQ_TX_IO_M1_CFG_3 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_3_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_3_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_3_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_3_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_3_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_3_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_3_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_3_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_3_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_3_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_3_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_3_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_3_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_3_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_3_ADR 32'h00000930
`define DDR_CA_DQ_TX_IO_M1_CFG_3_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_3_MSK 32'h00000FFF

// Word Address 0x00000934 : DDR_CA_DQ_TX_IO_M1_CFG_4 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_4_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_4_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_4_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_4_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_4_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_4_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_4_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_4_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_4_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_4_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_4_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_4_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_4_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_4_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_4_ADR 32'h00000934
`define DDR_CA_DQ_TX_IO_M1_CFG_4_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_4_MSK 32'h00000FFF

// Word Address 0x00000938 : DDR_CA_DQ_TX_IO_M1_CFG_5 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_5_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_5_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_5_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_5_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_5_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_5_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_5_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_5_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_5_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_5_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_5_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_5_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_5_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_5_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_5_ADR 32'h00000938
`define DDR_CA_DQ_TX_IO_M1_CFG_5_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_5_MSK 32'h00000FFF

// Word Address 0x0000093C : DDR_CA_DQ_TX_IO_M1_CFG_6 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_6_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_6_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_6_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_6_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_6_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_6_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_6_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_6_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_6_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_6_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_6_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_6_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_6_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_6_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_6_ADR 32'h0000093C
`define DDR_CA_DQ_TX_IO_M1_CFG_6_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_6_MSK 32'h00000FFF

// Word Address 0x00000940 : DDR_CA_DQ_TX_IO_M1_CFG_7 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_7_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_7_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_7_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_7_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_7_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_7_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_7_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_7_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_7_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_7_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_7_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_7_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_7_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_7_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_7_ADR 32'h00000940
`define DDR_CA_DQ_TX_IO_M1_CFG_7_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_7_MSK 32'h00000FFF

// Word Address 0x00000944 : DDR_CA_DQ_TX_IO_M1_CFG_8 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_8_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_8_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_8_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_8_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_8_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_8_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_8_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_8_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_8_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_8_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_8_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_8_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_8_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_8_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_8_ADR 32'h00000944
`define DDR_CA_DQ_TX_IO_M1_CFG_8_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_8_MSK 32'h00000FFF

// Word Address 0x00000948 : DDR_CA_DQ_TX_IO_M1_CFG_9 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_9_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_9_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_9_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_9_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_9_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_9_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_9_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_9_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_9_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_9_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_9_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_9_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_9_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_9_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_9_ADR 32'h00000948
`define DDR_CA_DQ_TX_IO_M1_CFG_9_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_9_MSK 32'h00000FFF

// Word Address 0x0000094C : DDR_CA_DQ_TX_IO_M1_CFG_10 (RW)
`define DDR_CA_DQ_TX_IO_M1_CFG_10_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQ_TX_IO_M1_CFG_10_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_10_OVRD_VAL_FIELD 3
`define DDR_CA_DQ_TX_IO_M1_CFG_10_OVRD_VAL_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_10_RESERVED_FIELD 4
`define DDR_CA_DQ_TX_IO_M1_CFG_10_RESERVED_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_10_RX_IMPD_FIELD 11:9
`define DDR_CA_DQ_TX_IO_M1_CFG_10_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_10_SW_OVR_FIELD 5
`define DDR_CA_DQ_TX_IO_M1_CFG_10_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQ_TX_IO_M1_CFG_10_TX_IMPD_FIELD 8:6
`define DDR_CA_DQ_TX_IO_M1_CFG_10_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQ_TX_IO_M1_CFG_10_RANGE 11:0
`define DDR_CA_DQ_TX_IO_M1_CFG_10_WIDTH 12
`define DDR_CA_DQ_TX_IO_M1_CFG_10_ADR 32'h0000094C
`define DDR_CA_DQ_TX_IO_M1_CFG_10_POR 32'h00000040
`define DDR_CA_DQ_TX_IO_M1_CFG_10_MSK 32'h00000FFF

// Word Address 0x00000950 : DDR_CA_DQS_RX_M0_CFG (RW)
`define DDR_CA_DQS_RX_M0_CFG_FGB_MODE_FIELD 7:4
`define DDR_CA_DQS_RX_M0_CFG_FGB_MODE_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_M0_CFG_PRE_FILTER_SEL_FIELD 13:12
`define DDR_CA_DQS_RX_M0_CFG_PRE_FILTER_SEL_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_M0_CFG_RGB_MODE_FIELD 2:0
`define DDR_CA_DQS_RX_M0_CFG_RGB_MODE_FIELD_WIDTH 3
`define DDR_CA_DQS_RX_M0_CFG_WCK_MODE_FIELD 8
`define DDR_CA_DQS_RX_M0_CFG_WCK_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_M0_CFG_RANGE 13:0
`define DDR_CA_DQS_RX_M0_CFG_WIDTH 14
`define DDR_CA_DQS_RX_M0_CFG_ADR 32'h00000950
`define DDR_CA_DQS_RX_M0_CFG_POR 32'h00000074
`define DDR_CA_DQS_RX_M0_CFG_MSK 32'h000031F7

// Word Address 0x00000954 : DDR_CA_DQS_RX_M1_CFG (RW)
`define DDR_CA_DQS_RX_M1_CFG_FGB_MODE_FIELD 7:4
`define DDR_CA_DQS_RX_M1_CFG_FGB_MODE_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_M1_CFG_PRE_FILTER_SEL_FIELD 13:12
`define DDR_CA_DQS_RX_M1_CFG_PRE_FILTER_SEL_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_M1_CFG_RGB_MODE_FIELD 2:0
`define DDR_CA_DQS_RX_M1_CFG_RGB_MODE_FIELD_WIDTH 3
`define DDR_CA_DQS_RX_M1_CFG_WCK_MODE_FIELD 8
`define DDR_CA_DQS_RX_M1_CFG_WCK_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_M1_CFG_RANGE 13:0
`define DDR_CA_DQS_RX_M1_CFG_WIDTH 14
`define DDR_CA_DQS_RX_M1_CFG_ADR 32'h00000954
`define DDR_CA_DQS_RX_M1_CFG_POR 32'h00000074
`define DDR_CA_DQS_RX_M1_CFG_MSK 32'h000031F7

// Word Address 0x00000958 : DDR_CA_DQS_RX_BSCAN_STA (R)
`define DDR_CA_DQS_RX_BSCAN_STA_VAL_FIELD 1:0
`define DDR_CA_DQS_RX_BSCAN_STA_VAL_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_BSCAN_STA_RANGE 1:0
`define DDR_CA_DQS_RX_BSCAN_STA_WIDTH 2
`define DDR_CA_DQS_RX_BSCAN_STA_ADR 32'h00000958
`define DDR_CA_DQS_RX_BSCAN_STA_POR 32'h00000000
`define DDR_CA_DQS_RX_BSCAN_STA_MSK 32'h00000003

// Word Address 0x0000095C : DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG (RW)
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_EN_FIELD 8
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_GEAR_FIELD 7:6
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_RANGE 8:0
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_WIDTH 9
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_ADR 32'h0000095C
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_POR 32'h00000100
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R0_CFG_MSK 32'h000001FF

// Word Address 0x00000960 : DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG (RW)
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_EN_FIELD 8
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_GEAR_FIELD 7:6
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_RANGE 8:0
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_WIDTH 9
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_ADR 32'h00000960
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_POR 32'h00000100
`define DDR_CA_DQS_RX_SDR_LPDE_M0_R1_CFG_MSK 32'h000001FF

// Word Address 0x00000964 : DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG (RW)
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_EN_FIELD 8
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_GEAR_FIELD 7:6
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_RANGE 8:0
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_WIDTH 9
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_ADR 32'h00000964
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_POR 32'h00000100
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R0_CFG_MSK 32'h000001FF

// Word Address 0x00000968 : DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG (RW)
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_EN_FIELD 8
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_GEAR_FIELD 7:6
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_RANGE 8:0
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_WIDTH 9
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_ADR 32'h00000968
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_POR 32'h00000100
`define DDR_CA_DQS_RX_SDR_LPDE_M1_R1_CFG_MSK 32'h000001FF

// Word Address 0x0000096C : DDR_CA_DQS_RX_REN_PI_M0_R0_CFG (RW)
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_ADR 32'h0000096C
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_REN_PI_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000970 : DDR_CA_DQS_RX_REN_PI_M0_R1_CFG (RW)
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_ADR 32'h00000970
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_REN_PI_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000974 : DDR_CA_DQS_RX_REN_PI_M1_R0_CFG (RW)
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_ADR 32'h00000974
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_REN_PI_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000978 : DDR_CA_DQS_RX_REN_PI_M1_R1_CFG (RW)
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_ADR 32'h00000978
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_REN_PI_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x0000097C : DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG (RW)
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_ADR 32'h0000097C
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RCS_PI_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000980 : DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG (RW)
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_ADR 32'h00000980
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RCS_PI_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000984 : DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG (RW)
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_ADR 32'h00000984
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RCS_PI_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000988 : DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG (RW)
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_ADR 32'h00000988
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RCS_PI_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x0000098C : DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_ADR 32'h0000098C
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000990 : DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_ADR 32'h00000990
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_0_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000994 : DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_ADR 32'h00000994
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000998 : DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_ADR 32'h00000998
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_0_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x0000099C : DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_ADR 32'h0000099C
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x000009A0 : DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_ADR 32'h000009A0
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_1_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x000009A4 : DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_ADR 32'h000009A4
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x000009A8 : DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG (RW)
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_ADR 32'h000009A8
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_RX_RDQS_PI_1_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x000009AC : DDR_CA_DQS_RX_PI_STA (R)
`define DDR_CA_DQS_RX_PI_STA_RCS_PI_PHASE_FIELD 1
`define DDR_CA_DQS_RX_PI_STA_RCS_PI_PHASE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_PI_STA_REN_PI_PHASE_FIELD 0
`define DDR_CA_DQS_RX_PI_STA_REN_PI_PHASE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_PI_STA_RANGE 1:0
`define DDR_CA_DQS_RX_PI_STA_WIDTH 2
`define DDR_CA_DQS_RX_PI_STA_ADR 32'h000009AC
`define DDR_CA_DQS_RX_PI_STA_POR 32'h00000000
`define DDR_CA_DQS_RX_PI_STA_MSK 32'h00000003

// Word Address 0x000009B0 : DDR_CA_DQS_RX_IO_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_DLY_CTRL_C_FIELD 7:0
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_DLY_CTRL_C_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_DLY_CTRL_T_FIELD 15:8
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_DLY_CTRL_T_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_RANGE 15:0
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_WIDTH 16
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_ADR 32'h000009B0
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_IO_M0_R0_CFG_0_MSK 32'h0000FFFF

// Word Address 0x000009B4 : DDR_CA_DQS_RX_IO_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_DLY_CTRL_C_FIELD 7:0
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_DLY_CTRL_C_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_DLY_CTRL_T_FIELD 15:8
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_DLY_CTRL_T_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_RANGE 15:0
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_WIDTH 16
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_ADR 32'h000009B4
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_IO_M0_R1_CFG_0_MSK 32'h0000FFFF

// Word Address 0x000009B8 : DDR_CA_DQS_RX_IO_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_DLY_CTRL_C_FIELD 7:0
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_DLY_CTRL_C_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_DLY_CTRL_T_FIELD 15:8
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_DLY_CTRL_T_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_RANGE 15:0
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_WIDTH 16
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_ADR 32'h000009B8
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_IO_M1_R0_CFG_0_MSK 32'h0000FFFF

// Word Address 0x000009BC : DDR_CA_DQS_RX_IO_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_DLY_CTRL_C_FIELD 7:0
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_DLY_CTRL_C_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_DLY_CTRL_T_FIELD 15:8
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_DLY_CTRL_T_FIELD_WIDTH 8
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_RANGE 15:0
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_WIDTH 16
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_ADR 32'h000009BC
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_IO_M1_R1_CFG_0_MSK 32'h0000FFFF

// Word Address 0x000009C0 : DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG (RW)
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_N_C_FIELD 11:8
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_N_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_N_T_FIELD 15:12
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_N_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_P_C_FIELD 3:0
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_P_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_P_T_FIELD 7:4
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_CAL_P_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_DCPATH_EN_FIELD 19
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_DCPATH_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_EN_FIELD 20
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_FB_EN_FIELD 18:16
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_FB_EN_FIELD_WIDTH 3
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_RXCAL_EN_FIELD 21
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_RXCAL_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_SE_MODE_FIELD 22
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_SW_OVR_FIELD 23
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_RANGE 23:0
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_WIDTH 24
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_ADR 32'h000009C0
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_POR 32'h004A7777
`define DDR_CA_DQS_RX_IO_CMN_M0_R0_CFG_MSK 32'h00FFFFFF

// Word Address 0x000009C4 : DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG (RW)
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_N_C_FIELD 11:8
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_N_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_N_T_FIELD 15:12
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_N_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_P_C_FIELD 3:0
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_P_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_P_T_FIELD 7:4
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_CAL_P_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_DCPATH_EN_FIELD 19
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_DCPATH_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_EN_FIELD 20
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_FB_EN_FIELD 18:16
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_FB_EN_FIELD_WIDTH 3
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_RXCAL_EN_FIELD 21
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_RXCAL_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_SE_MODE_FIELD 22
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_SW_OVR_FIELD 23
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_RANGE 23:0
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_WIDTH 24
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_ADR 32'h000009C4
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_POR 32'h004A7777
`define DDR_CA_DQS_RX_IO_CMN_M0_R1_CFG_MSK 32'h00FFFFFF

// Word Address 0x000009C8 : DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG (RW)
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_N_C_FIELD 11:8
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_N_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_N_T_FIELD 15:12
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_N_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_P_C_FIELD 3:0
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_P_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_P_T_FIELD 7:4
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_CAL_P_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_DCPATH_EN_FIELD 19
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_DCPATH_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_EN_FIELD 20
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_FB_EN_FIELD 18:16
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_FB_EN_FIELD_WIDTH 3
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_RXCAL_EN_FIELD 21
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_RXCAL_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_SE_MODE_FIELD 22
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_SW_OVR_FIELD 23
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_RANGE 23:0
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_WIDTH 24
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_ADR 32'h000009C8
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_POR 32'h004A7777
`define DDR_CA_DQS_RX_IO_CMN_M1_R0_CFG_MSK 32'h00FFFFFF

// Word Address 0x000009CC : DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG (RW)
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_N_C_FIELD 11:8
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_N_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_N_T_FIELD 15:12
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_N_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_P_C_FIELD 3:0
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_P_C_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_P_T_FIELD 7:4
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_CAL_P_T_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_DCPATH_EN_FIELD 19
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_DCPATH_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_EN_FIELD 20
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_FB_EN_FIELD 18:16
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_FB_EN_FIELD_WIDTH 3
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_RXCAL_EN_FIELD 21
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_RXCAL_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_SE_MODE_FIELD 22
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_SW_OVR_FIELD 23
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_RANGE 23:0
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_WIDTH 24
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_ADR 32'h000009CC
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_POR 32'h004A7777
`define DDR_CA_DQS_RX_IO_CMN_M1_R1_CFG_MSK 32'h00FFFFFF

// Word Address 0x000009D0 : DDR_CA_DQS_RX_IO_STA (R)
`define DDR_CA_DQS_RX_IO_STA_CORE_IG_FIELD 31:0
`define DDR_CA_DQS_RX_IO_STA_CORE_IG_FIELD_WIDTH 32
`define DDR_CA_DQS_RX_IO_STA_RANGE 31:0
`define DDR_CA_DQS_RX_IO_STA_WIDTH 32
`define DDR_CA_DQS_RX_IO_STA_ADR 32'h000009D0
`define DDR_CA_DQS_RX_IO_STA_POR 32'h00000000
`define DDR_CA_DQS_RX_IO_STA_MSK 32'hFFFFFFFF

// Word Address 0x000009D4 : DDR_CA_DQS_RX_SA_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_RANGE 19:0
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_WIDTH 20
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_ADR 32'h000009D4
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_SA_M0_R0_CFG_0_MSK 32'h000FFFFF

// Word Address 0x000009D8 : DDR_CA_DQS_RX_SA_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_RANGE 19:0
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_WIDTH 20
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_ADR 32'h000009D8
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_SA_M0_R1_CFG_0_MSK 32'h000FFFFF

// Word Address 0x000009DC : DDR_CA_DQS_RX_SA_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_RANGE 19:0
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_WIDTH 20
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_ADR 32'h000009DC
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_SA_M1_R0_CFG_0_MSK 32'h000FFFFF

// Word Address 0x000009E0 : DDR_CA_DQS_RX_SA_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_0_FIELD 3:0
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_0_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_180_FIELD 11:8
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_180_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_270_FIELD 15:12
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_270_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_90_FIELD 7:4
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_CODE_90_FIELD_WIDTH 4
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_0_FIELD 16
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_0_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_180_FIELD 18
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_180_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_270_FIELD 19
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_270_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_90_FIELD 17
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_CAL_DIR_90_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_RANGE 19:0
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_WIDTH 20
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_ADR 32'h000009E0
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_RX_SA_M1_R1_CFG_0_MSK 32'h000FFFFF

// Word Address 0x000009E4 : DDR_CA_DQS_RX_SA_CMN_CFG (RW)
`define DDR_CA_DQS_RX_SA_CMN_CFG_CAL_EN_0_180_FIELD 1
`define DDR_CA_DQS_RX_SA_CMN_CFG_CAL_EN_0_180_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_CMN_CFG_CAL_EN_90_270_FIELD 3
`define DDR_CA_DQS_RX_SA_CMN_CFG_CAL_EN_90_270_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_CMN_CFG_OVR_EN_0_180_FIELD 0
`define DDR_CA_DQS_RX_SA_CMN_CFG_OVR_EN_0_180_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_CMN_CFG_OVR_EN_90_270_FIELD 2
`define DDR_CA_DQS_RX_SA_CMN_CFG_OVR_EN_90_270_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_CMN_CFG_SW_OVR_FIELD 4
`define DDR_CA_DQS_RX_SA_CMN_CFG_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_RX_SA_CMN_CFG_RANGE 4:0
`define DDR_CA_DQS_RX_SA_CMN_CFG_WIDTH 5
`define DDR_CA_DQS_RX_SA_CMN_CFG_ADR 32'h000009E4
`define DDR_CA_DQS_RX_SA_CMN_CFG_POR 32'h00000005
`define DDR_CA_DQS_RX_SA_CMN_CFG_MSK 32'h0000001F

// Word Address 0x000009E8 : DDR_CA_DQS_TX_M0_CFG (RW)
`define DDR_CA_DQS_TX_M0_CFG_CK2WCK_RATIO_FIELD 9:8
`define DDR_CA_DQS_TX_M0_CFG_CK2WCK_RATIO_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_M0_CFG_TGB_MODE_FIELD 2:0
`define DDR_CA_DQS_TX_M0_CFG_TGB_MODE_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_M0_CFG_WGB_MODE_FIELD 7:4
`define DDR_CA_DQS_TX_M0_CFG_WGB_MODE_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_M0_CFG_RANGE 9:0
`define DDR_CA_DQS_TX_M0_CFG_WIDTH 10
`define DDR_CA_DQS_TX_M0_CFG_ADR 32'h000009E8
`define DDR_CA_DQS_TX_M0_CFG_POR 32'h00000087
`define DDR_CA_DQS_TX_M0_CFG_MSK 32'h000003F7

// Word Address 0x000009EC : DDR_CA_DQS_TX_M1_CFG (RW)
`define DDR_CA_DQS_TX_M1_CFG_CK2WCK_RATIO_FIELD 9:8
`define DDR_CA_DQS_TX_M1_CFG_CK2WCK_RATIO_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_M1_CFG_TGB_MODE_FIELD 2:0
`define DDR_CA_DQS_TX_M1_CFG_TGB_MODE_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_M1_CFG_WGB_MODE_FIELD 7:4
`define DDR_CA_DQS_TX_M1_CFG_WGB_MODE_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_M1_CFG_RANGE 9:0
`define DDR_CA_DQS_TX_M1_CFG_WIDTH 10
`define DDR_CA_DQS_TX_M1_CFG_ADR 32'h000009EC
`define DDR_CA_DQS_TX_M1_CFG_POR 32'h00000087
`define DDR_CA_DQS_TX_M1_CFG_MSK 32'h000003F7

// Word Address 0x000009F0 : DDR_CA_DQS_TX_BSCAN_CTRL_CFG (RW)
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_IE_FIELD 0
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_IE_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_OE_FIELD 1
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_OE_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_RANGE 1:0
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_WIDTH 2
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_ADR 32'h000009F0
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_POR 32'h00000000
`define DDR_CA_DQS_TX_BSCAN_CTRL_CFG_MSK 32'h00000003

// Word Address 0x000009F4 : DDR_CA_DQS_TX_BSCAN_CFG (RW)
`define DDR_CA_DQS_TX_BSCAN_CFG_VAL_FIELD 1:0
`define DDR_CA_DQS_TX_BSCAN_CFG_VAL_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_BSCAN_CFG_RANGE 1:0
`define DDR_CA_DQS_TX_BSCAN_CFG_WIDTH 2
`define DDR_CA_DQS_TX_BSCAN_CFG_ADR 32'h000009F4
`define DDR_CA_DQS_TX_BSCAN_CFG_POR 32'h00000000
`define DDR_CA_DQS_TX_BSCAN_CFG_MSK 32'h00000003

// Word Address 0x000009F8 : DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0 (RW)
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_RANGE 5:0
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_WIDTH 6
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_ADR 32'h000009F8
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_POR 32'h00000001
`define DDR_CA_DQS_TX_EGRESS_ANA_M0_CFG_0_MSK 32'h0000003F

// Word Address 0x000009FC : DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0 (RW)
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_EGRESS_MODE_FIELD 5:0
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_EGRESS_MODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_RANGE 5:0
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_WIDTH 6
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_ADR 32'h000009FC
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_POR 32'h00000001
`define DDR_CA_DQS_TX_EGRESS_ANA_M1_CFG_0_MSK 32'h0000003F

// Word Address 0x00000A00 : DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0 (RW)
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_RANGE 6:0
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_WIDTH 7
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_ADR 32'h00000A00
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_POR 32'h00000002
`define DDR_CA_DQS_TX_EGRESS_DIG_M0_CFG_0_MSK 32'h0000007F

// Word Address 0x00000A04 : DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0 (RW)
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_EGRESS_MODE_FIELD 6:0
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_EGRESS_MODE_FIELD_WIDTH 7
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_RANGE 6:0
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_WIDTH 7
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_ADR 32'h00000A04
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_POR 32'h00000002
`define DDR_CA_DQS_TX_EGRESS_DIG_M1_CFG_0_MSK 32'h0000007F

// Word Address 0x00000A08 : DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_ADR 32'h00000A08
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_ODR_PI_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A0C : DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_ADR 32'h00000A0C
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_ODR_PI_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A10 : DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_ADR 32'h00000A10
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_ODR_PI_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A14 : DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_ADR 32'h00000A14
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_ODR_PI_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A18 : DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_ADR 32'h00000A18
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A1C : DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_ADR 32'h00000A1C
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_0_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A20 : DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_ADR 32'h00000A20
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A24 : DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_ADR 32'h00000A24
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_0_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A28 : DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_ADR 32'h00000A28
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A2C : DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_ADR 32'h00000A2C
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_1_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A30 : DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_ADR 32'h00000A30
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A34 : DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_ADR 32'h00000A34
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_QDR_PI_1_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A38 : DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_ADR 32'h00000A38
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A3C : DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_ADR 32'h00000A3C
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_0_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A40 : DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_ADR 32'h00000A40
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A44 : DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_ADR 32'h00000A44
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_0_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A48 : DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_ADR 32'h00000A48
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A4C : DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_ADR 32'h00000A4C
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_1_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A50 : DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_ADR 32'h00000A50
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A54 : DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_ADR 32'h00000A54
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DDR_PI_1_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A58 : DDR_CA_DQS_TX_PI_RT_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_ADR 32'h00000A58
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_PI_RT_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A5C : DDR_CA_DQS_TX_PI_RT_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_ADR 32'h00000A5C
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_PI_RT_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A60 : DDR_CA_DQS_TX_PI_RT_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_ADR 32'h00000A60
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_PI_RT_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A64 : DDR_CA_DQS_TX_PI_RT_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_CODE_FIELD 5:0
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_CODE_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_ADR 32'h00000A64
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_PI_RT_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A68 : DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_ADR 32'h00000A68
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_SDR_PI_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A6C : DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_ADR 32'h00000A6C
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_SDR_PI_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A70 : DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_ADR 32'h00000A70
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_SDR_PI_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A74 : DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_ADR 32'h00000A74
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_SDR_PI_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A78 : DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_ADR 32'h00000A78
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DFI_PI_M0_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A7C : DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_ADR 32'h00000A7C
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DFI_PI_M0_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A80 : DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_ADR 32'h00000A80
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DFI_PI_M1_R0_CFG_MSK 32'h00007FFF

// Word Address 0x00000A84 : DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_EN_FIELD 14
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_GEAR_FIELD 9:6
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_GEAR_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_RSVD_FIELD 5:0
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_RSVD_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_XCPL_FIELD 13:10
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_XCPL_FIELD_WIDTH 4
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_RANGE 14:0
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_WIDTH 15
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_ADR 32'h00000A84
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_POR 32'h00000040
`define DDR_CA_DQS_TX_DFI_PI_M1_R1_CFG_MSK 32'h00007FFF

// Word Address 0x00000A88 : DDR_CA_DQS_TX_RT_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_PIPE_EN_FIELD 0:0
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_RANGE 0:0
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_WIDTH 1
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_ADR 32'h00000A88
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_POR 32'h00000000
`define DDR_CA_DQS_TX_RT_M0_R0_CFG_MSK 32'h00000001

// Word Address 0x00000A8C : DDR_CA_DQS_TX_RT_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_PIPE_EN_FIELD 0:0
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_RANGE 0:0
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_WIDTH 1
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_ADR 32'h00000A8C
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_POR 32'h00000000
`define DDR_CA_DQS_TX_RT_M0_R1_CFG_MSK 32'h00000001

// Word Address 0x00000A90 : DDR_CA_DQS_TX_RT_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_PIPE_EN_FIELD 0:0
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_RANGE 0:0
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_WIDTH 1
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_ADR 32'h00000A90
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_POR 32'h00000000
`define DDR_CA_DQS_TX_RT_M1_R0_CFG_MSK 32'h00000001

// Word Address 0x00000A94 : DDR_CA_DQS_TX_RT_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_PIPE_EN_FIELD 0:0
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_PIPE_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_RANGE 0:0
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_WIDTH 1
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_ADR 32'h00000A94
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_POR 32'h00000000
`define DDR_CA_DQS_TX_RT_M1_R1_CFG_MSK 32'h00000001

// Word Address 0x00000A98 : DDR_CA_DQS_TX_SDR_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_RANGE 7:0
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_WIDTH 8
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_ADR 32'h00000A98
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_M0_R0_CFG_0_MSK 32'h000000FF

// Word Address 0x00000A9C : DDR_CA_DQS_TX_SDR_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_RANGE 7:0
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_WIDTH 8
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_ADR 32'h00000A9C
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_M0_R1_CFG_0_MSK 32'h000000FF

// Word Address 0x00000AA0 : DDR_CA_DQS_TX_SDR_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_RANGE 7:0
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_WIDTH 8
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_ADR 32'h00000AA0
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_M1_R0_CFG_0_MSK 32'h000000FF

// Word Address 0x00000AA4 : DDR_CA_DQS_TX_SDR_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P4_FIELD 4
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P4_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P5_FIELD 5
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P5_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P6_FIELD 6
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P6_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P7_FIELD 7
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_PIPE_EN_P7_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_RANGE 7:0
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_WIDTH 8
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_ADR 32'h00000AA4
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_M1_R1_CFG_0_MSK 32'h000000FF

// Word Address 0x00000AA8 : DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_RANGE 30:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_WIDTH 31
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_ADR 32'h00000AA8
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R0_CFG_0_MSK 32'h77777777

// Word Address 0x00000AAC : DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_RANGE 30:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_WIDTH 31
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_ADR 32'h00000AAC
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_X_SEL_M0_R1_CFG_0_MSK 32'h77777777

// Word Address 0x00000AB0 : DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_RANGE 30:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_WIDTH 31
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_ADR 32'h00000AB0
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R0_CFG_0_MSK 32'h77777777

// Word Address 0x00000AB4 : DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD 2:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD 6:4
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD 10:8
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD 14:12
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P4_FIELD 18:16
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P4_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P5_FIELD 22:20
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P5_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P6_FIELD 26:24
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P6_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P7_FIELD 30:28
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_X_SEL_P7_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_RANGE 30:0
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_WIDTH 31
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_ADR 32'h00000AB4
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_X_SEL_M1_R1_CFG_0_MSK 32'h77777777

// Word Address 0x00000AB8 : DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_RANGE 29:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_WIDTH 30
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_ADR 32'h00000AB8
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0_MSK 32'h33333333

// Word Address 0x00000ABC : DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_RANGE 29:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_WIDTH 30
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_ADR 32'h00000ABC
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0_MSK 32'h33333333

// Word Address 0x00000AC0 : DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_RANGE 29:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_WIDTH 30
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_ADR 32'h00000AC0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0_MSK 32'h33333333

// Word Address 0x00000AC4 : DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P0_FIELD 1:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P1_FIELD 5:4
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P2_FIELD 9:8
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P3_FIELD 13:12
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P4_FIELD 17:16
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P4_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P5_FIELD 21:20
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P5_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P6_FIELD 25:24
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P6_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P7_FIELD 29:28
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_DLY_P7_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_RANGE 29:0
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_WIDTH 30
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_ADR 32'h00000AC4
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0_MSK 32'h33333333

// Word Address 0x00000AC8 : DDR_CA_DQS_TX_DDR_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_RANGE 3:0
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_WIDTH 4
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_ADR 32'h00000AC8
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_M0_R0_CFG_0_MSK 32'h0000000F

// Word Address 0x00000ACC : DDR_CA_DQS_TX_DDR_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_RANGE 3:0
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_WIDTH 4
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_ADR 32'h00000ACC
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_M0_R1_CFG_0_MSK 32'h0000000F

// Word Address 0x00000AD0 : DDR_CA_DQS_TX_DDR_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_RANGE 3:0
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_WIDTH 4
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_ADR 32'h00000AD0
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_M1_R0_CFG_0_MSK 32'h0000000F

// Word Address 0x00000AD4 : DDR_CA_DQS_TX_DDR_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD 2
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P2_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD 3
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_PIPE_EN_P3_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_RANGE 3:0
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_WIDTH 4
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_ADR 32'h00000AD4
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_M1_R1_CFG_0_MSK 32'h0000000F

// Word Address 0x00000AD8 : DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_RANGE 13:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_WIDTH 14
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_ADR 32'h00000AD8
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R0_CFG_0_MSK 32'h00003333

// Word Address 0x00000ADC : DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_RANGE 13:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_WIDTH 14
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_ADR 32'h00000ADC
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_X_SEL_M0_R1_CFG_0_MSK 32'h00003333

// Word Address 0x00000AE0 : DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_RANGE 13:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_WIDTH 14
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_ADR 32'h00000AE0
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R0_CFG_0_MSK 32'h00003333

// Word Address 0x00000AE4 : DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD 1:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD 5:4
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD 9:8
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P2_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD 13:12
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_X_SEL_P3_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_RANGE 13:0
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_WIDTH 14
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_ADR 32'h00000AE4
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_DDR_X_SEL_M1_R1_CFG_0_MSK 32'h00003333

// Word Address 0x00000AE8 : DDR_CA_DQS_TX_QDR_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_RANGE 1:0
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_WIDTH 2
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_ADR 32'h00000AE8
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_M0_R0_CFG_0_MSK 32'h00000003

// Word Address 0x00000AEC : DDR_CA_DQS_TX_QDR_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_RANGE 1:0
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_WIDTH 2
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_ADR 32'h00000AEC
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_M0_R1_CFG_0_MSK 32'h00000003

// Word Address 0x00000AF0 : DDR_CA_DQS_TX_QDR_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_RANGE 1:0
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_WIDTH 2
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_ADR 32'h00000AF0
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_M1_R0_CFG_0_MSK 32'h00000003

// Word Address 0x00000AF4 : DDR_CA_DQS_TX_QDR_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_PIPE_EN_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD 1
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_PIPE_EN_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_RANGE 1:0
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_WIDTH 2
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_ADR 32'h00000AF4
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_M1_R1_CFG_0_MSK 32'h00000003

// Word Address 0x00000AF8 : DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_RANGE 4:0
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_WIDTH 5
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_ADR 32'h00000AF8
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R0_CFG_0_MSK 32'h00000011

// Word Address 0x00000AFC : DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_RANGE 4:0
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_WIDTH 5
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_ADR 32'h00000AFC
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_X_SEL_M0_R1_CFG_0_MSK 32'h00000011

// Word Address 0x00000B00 : DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_RANGE 4:0
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_WIDTH 5
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_ADR 32'h00000B00
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R0_CFG_0_MSK 32'h00000011

// Word Address 0x00000B04 : DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD 0
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P0_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD 4
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_X_SEL_P1_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_RANGE 4:0
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_WIDTH 5
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_ADR 32'h00000B04
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_POR 32'h00000000
`define DDR_CA_DQS_TX_QDR_X_SEL_M1_R1_CFG_0_MSK 32'h00000011

// Word Address 0x00000B08 : DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_EN_FIELD 8
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_RANGE 8:0
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_WIDTH 9
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_ADR 32'h00000B08
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_POR 32'h00000100
`define DDR_CA_DQS_TX_LPDE_M0_R0_CFG_0_MSK 32'h000001FF

// Word Address 0x00000B0C : DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_EN_FIELD 8
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_RANGE 8:0
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_WIDTH 9
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_ADR 32'h00000B0C
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_POR 32'h00000100
`define DDR_CA_DQS_TX_LPDE_M0_R1_CFG_0_MSK 32'h000001FF

// Word Address 0x00000B10 : DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0 (RW)
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_EN_FIELD 8
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_RANGE 8:0
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_WIDTH 9
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_ADR 32'h00000B10
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_POR 32'h00000100
`define DDR_CA_DQS_TX_LPDE_M1_R0_CFG_0_MSK 32'h000001FF

// Word Address 0x00000B14 : DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0 (RW)
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_CTRL_BIN_FIELD 5:0
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_CTRL_BIN_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_EN_FIELD 8
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_GEAR_FIELD 7:6
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_GEAR_FIELD_WIDTH 2
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_RANGE 8:0
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_WIDTH 9
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_ADR 32'h00000B14
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_POR 32'h00000100
`define DDR_CA_DQS_TX_LPDE_M1_R1_CFG_0_MSK 32'h000001FF

// Word Address 0x00000B18 : DDR_CA_DQS_TX_IO_M0_CFG_0 (RW)
`define DDR_CA_DQS_TX_IO_M0_CFG_0_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQS_TX_IO_M0_CFG_0_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_IO_M0_CFG_0_OVRD_VAL_C_FIELD 3
`define DDR_CA_DQS_TX_IO_M0_CFG_0_OVRD_VAL_C_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_M0_CFG_0_OVRD_VAL_T_FIELD 4
`define DDR_CA_DQS_TX_IO_M0_CFG_0_OVRD_VAL_T_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_M0_CFG_0_RX_IMPD_FIELD 11:9
`define DDR_CA_DQS_TX_IO_M0_CFG_0_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_IO_M0_CFG_0_SW_OVR_FIELD 5
`define DDR_CA_DQS_TX_IO_M0_CFG_0_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_M0_CFG_0_TX_IMPD_FIELD 8:6
`define DDR_CA_DQS_TX_IO_M0_CFG_0_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_IO_M0_CFG_0_RANGE 11:0
`define DDR_CA_DQS_TX_IO_M0_CFG_0_WIDTH 12
`define DDR_CA_DQS_TX_IO_M0_CFG_0_ADR 32'h00000B18
`define DDR_CA_DQS_TX_IO_M0_CFG_0_POR 32'h00000041
`define DDR_CA_DQS_TX_IO_M0_CFG_0_MSK 32'h00000FFF

// Word Address 0x00000B1C : DDR_CA_DQS_TX_IO_M1_CFG_0 (RW)
`define DDR_CA_DQS_TX_IO_M1_CFG_0_OVRD_SEL_FIELD 2:0
`define DDR_CA_DQS_TX_IO_M1_CFG_0_OVRD_SEL_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_IO_M1_CFG_0_OVRD_VAL_C_FIELD 3
`define DDR_CA_DQS_TX_IO_M1_CFG_0_OVRD_VAL_C_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_M1_CFG_0_OVRD_VAL_T_FIELD 4
`define DDR_CA_DQS_TX_IO_M1_CFG_0_OVRD_VAL_T_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_M1_CFG_0_RX_IMPD_FIELD 11:9
`define DDR_CA_DQS_TX_IO_M1_CFG_0_RX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_IO_M1_CFG_0_SW_OVR_FIELD 5
`define DDR_CA_DQS_TX_IO_M1_CFG_0_SW_OVR_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_M1_CFG_0_TX_IMPD_FIELD 8:6
`define DDR_CA_DQS_TX_IO_M1_CFG_0_TX_IMPD_FIELD_WIDTH 3
`define DDR_CA_DQS_TX_IO_M1_CFG_0_RANGE 11:0
`define DDR_CA_DQS_TX_IO_M1_CFG_0_WIDTH 12
`define DDR_CA_DQS_TX_IO_M1_CFG_0_ADR 32'h00000B1C
`define DDR_CA_DQS_TX_IO_M1_CFG_0_POR 32'h00000041
`define DDR_CA_DQS_TX_IO_M1_CFG_0_MSK 32'h00000FFF

// Word Address 0x00000B20 : DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG (RW)
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_BS_EN_FIELD 11
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_BS_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_LPBK_EN_FIELD 12
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_LPBK_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_NCAL_FIELD 4:0
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_NCAL_FIELD_WIDTH 5
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_PCAL_FIELD 10:5
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_PCAL_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_SE_MODE_FIELD 13
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_RANGE 13:0
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_WIDTH 14
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_ADR 32'h00000B20
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_POR 32'h00000001
`define DDR_CA_DQS_TX_IO_CMN_M0_R0_CFG_MSK 32'h00003FFF

// Word Address 0x00000B24 : DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG (RW)
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_BS_EN_FIELD 11
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_BS_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_LPBK_EN_FIELD 12
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_LPBK_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_NCAL_FIELD 4:0
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_NCAL_FIELD_WIDTH 5
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_PCAL_FIELD 10:5
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_PCAL_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_SE_MODE_FIELD 13
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_RANGE 13:0
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_WIDTH 14
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_ADR 32'h00000B24
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_POR 32'h00000001
`define DDR_CA_DQS_TX_IO_CMN_M0_R1_CFG_MSK 32'h00003FFF

// Word Address 0x00000B28 : DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG (RW)
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_BS_EN_FIELD 11
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_BS_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_LPBK_EN_FIELD 12
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_LPBK_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_NCAL_FIELD 4:0
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_NCAL_FIELD_WIDTH 5
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_PCAL_FIELD 10:5
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_PCAL_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_SE_MODE_FIELD 13
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_RANGE 13:0
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_WIDTH 14
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_ADR 32'h00000B28
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_POR 32'h00000001
`define DDR_CA_DQS_TX_IO_CMN_M1_R0_CFG_MSK 32'h00003FFF

// Word Address 0x00000B2C : DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG (RW)
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_BS_EN_FIELD 11
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_BS_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_LPBK_EN_FIELD 12
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_LPBK_EN_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_NCAL_FIELD 4:0
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_NCAL_FIELD_WIDTH 5
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_PCAL_FIELD 10:5
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_PCAL_FIELD_WIDTH 6
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_SE_MODE_FIELD 13
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_SE_MODE_FIELD_WIDTH 1
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_RANGE 13:0
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_WIDTH 14
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_ADR 32'h00000B2C
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_POR 32'h00000001
`define DDR_CA_DQS_TX_IO_CMN_M1_R1_CFG_MSK 32'h00003FFF
