/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 13323
// Design library name: wphy_gf12lp_lp4x5_sim_lib
// Design cell name: wphy_lp4x5_cmn_clks_svt_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wavshared_gf12lp_dig_lib, Cell - wphy_lp4x5_cmn_clks_svt_FFRES_DEMET_D1_GL16_RVT,
//View - schematic
// LAST TIME SAVED: Nov 10 10:24:09 2020
// NETLIST TIME: Dec  7 22:24:41 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_FFRES_DEMET_D1_GL16_RVT (q, vdd, vss, clk, clkb, d, rst, rstb, 
    tiehi, tielo);

output  q;

inout  vdd, vss;

input  clk, clkb, d, rst, rstb, tiehi, tielo;


wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT FF0 ( .tielo(tielo), .tiehi(tiehi), .rst(rst), 
    .vss(vss), .vdd(vdd), .rstb(rstb), .d(d), .clkb(clkb), .clk(clk), 
    .q(q_mid));

wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT FF1 ( .tielo(tielo), .tiehi(tiehi), .rst(rst), 
    .vss(vss), .vdd(vdd), .rstb(rstb), .d(q_mid), .clkb(clkb), 
    .clk(clk), .q(q));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt, View -
//schematic
// LAST TIME SAVED: Sep 17 20:49:50 2020
// NETLIST TIME: Dec  7 22:24:41 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt (o_clk, o_clk_b, vdd, vss, ena, i_clk, 
    i_clk_b);

output  o_clk, o_clk_b;

inout  vdd, vss;

input  ena, i_clk, i_clk_b;


wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT0 ( .out(ckb), .en(en), .enb(enb), .vss(vss), 
    .in(i_clk), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT1 ( .out(ckbb), .en(en), .enb(enb), .vss(vss), 
    .in(i_clk_b), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_TIELO_D2_GL16_RVT I1 ( .tielo(tielo), .vss(vss), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_PU_D1_GL16_RVT PU0 ( .vdd(vdd), .en(en), .y(ckb));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV3 ( .in(ena), .vss(vss), .out(net012), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1_1 ( .in(ckb), .vss(vss), .out(o_clk), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1_0 ( .in(ckb), .vss(vss), .out(o_clk), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(enb), .vss(vss), .out(en), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2_1 ( .in(ckbb), .vss(vss), .out(o_clk_b), 
    .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2_0 ( .in(ckbb), .vss(vss), .out(o_clk_b), 
    .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_PD_D1_GL16_RVT PD0 ( .vss(vss), .enb(enb), .y(ckbb));

wphy_lp4x5_cmn_clks_svt_TIEHI_D2_GL16_RVT I0 ( .tiehi(tiehi), .vss(vss), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_LAT_D1_GL16_RVT LA0 ( .tielo(tielo), .vss(vss), .vdd(vdd), 
    .tiehi(tiehi), .d(net012), .clkb(i_clk_b), .clk(i_clk), .q(enb));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_lp4x5_cmn_clks_svt_wphy_clk_div2_4g_core_svt,
//View - schematic
// LAST TIME SAVED: Sep 17 20:50:32 2020
// NETLIST TIME: Dec  7 22:24:41 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_wphy_clk_div2_4g_core_svt (o_clk0, o_clk90, o_clk180, o_clk270, 
    vdda, vss, i_byp, i_clk0, i_clk180, i_rst);

output  o_clk0, o_clk90, o_clk180, o_clk270;

inout  vdda, vss;

input  i_byp, i_clk0, i_clk180, i_rst;


wphy_lp4x5_cmn_clks_svt_TIELO_D2_GL16_RVT I6 ( .tielo(tielo), .vss(vss), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT NOR0 ( .tielo(tielo), .tiehi(tiehi), .y(rst_or_byp_n), 
    .vss(vss), .vdd(vdda), .b(i_byp), .a(i_rst));

wphy_lp4x5_cmn_clks_svt_TIEHI_D2_GL16_RVT I5 ( .tiehi(tiehi), .vss(vss), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV16 ( .in(x90), .vss(vss), .out(x270), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV19 ( .in(net021), .vss(vss), .out(o_clk0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV18 ( .in(net029), .vss(vss), .out(o_clk270), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV17 ( .in(net028), .vss(vss), .out(o_clk90), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV14 ( .in(x180), .vss(vss), .out(x0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV20 ( .in(net030), .vss(vss), .out(o_clk180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1 ( .in(bypb), .vss(vss), .out(bypa), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(i_byp), .vss(vss), .out(bypb), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV15 ( .in(net020), .vss(vss), .out(x90), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2 ( .in(net015), .vss(vss), .out(x180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV9 ( .in(rst_or_byp_n), .vss(vss), .out(rst_or_byp), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT I3 ( .out(net028), .en(bypa), .enb(bypb), .vss(vss), 
    .in(i_clk180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT3 ( .out(net021), .en(bypa), .enb(bypb), 
    .vss(vss), .in(i_clk0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT2 ( .out(net021), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT8 ( .out(net028), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x90), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT1 ( .out(net030), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT7 ( .out(net029), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x270), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT0 ( .out(net030), .en(bypa), .enb(bypb), 
    .vss(vss), .in(i_clk180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT I4 ( .out(net029), .en(bypa), .enb(bypb), .vss(vss), 
    .in(i_clk0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LAT0 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdda), .rstb(rst_or_byp_n), .d(net020), .clkb(i_clk0), 
    .clk(i_clk180), .q(net015));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LAT1 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdda), .rstb(rst_or_byp_n), .d(x180), .clkb(i_clk180), 
    .clk(i_clk0), .q(net020));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt, View -
//schematic
// LAST TIME SAVED: Dec  2 23:53:28 2020
// NETLIST TIME: Dec  7 22:24:41 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt (clka_sel, clkb_sel, o_clk0, o_clk180, vdda, vss, 
    clk_sel, ena, i_clka0, i_clka180, i_clkb0, i_clkb180);

output  clka_sel, clkb_sel, o_clk0, o_clk180;

inout  vdda, vss;

input  clk_sel, ena, i_clka0, i_clka180, i_clkb0, i_clkb180;


wphy_lp4x5_cmn_clks_svt_TIEHI_D2_GL16_RVT I2 ( .tiehi(tiehi), .vss(vss), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA1 ( .tielo(tielo), .set(enb), .vss(vss), 
    .vdd(vdda), .tiehi(tiehi), .d(net6), .clkb(clka180), .clk(clka0), 
    .q(net023));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA4 ( .tielo(tielo), .set(enb), .vss(vss), 
    .vdd(vdda), .tiehi(tiehi), .d(net3), .clkb(clkb180), .clk(clkb0), 
    .q(net022));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA2 ( .tielo(tielo), .set(enb), .vss(vss), 
    .vdd(vdda), .tiehi(tiehi), .d(net023), .clkb(clka0), .clk(clka180), 
    .q(net5));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA3 ( .tielo(tielo), .set(enb), .vss(vss), 
    .vdd(vdda), .tiehi(tiehi), .d(net022), .clkb(clkb0), .clk(clkb180), 
    .q(net2));

wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT LA02 ( .prst(enb), .prstb(en), .tielo(tielo), 
    .vss(vss), .vdd(vdda), .tiehi(tiehi), .d(y), .clkb(clkb180), 
    .clk(clkb0), .q(net3));

wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT LA01 ( .prst(enb), .prstb(en), .tielo(tielo), 
    .vss(vss), .vdd(vdda), .tiehi(tiehi), .d(net4), .clkb(clka180), 
    .clk(clka0), .q(net6));

wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT NAND2 ( .tielo(tielo), .vdd(vdda), .y(pu_en), 
    .vss(vss), .tiehi(tiehi), .b(enb_b), .a(enb_a));

wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT NAND1 ( .tielo(tielo), .vdd(vdda), .y(y), .vss(vss), 
    .tiehi(tiehi), .b(net5), .a(sel_clkb));

wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT NAND0 ( .tielo(tielo), .vdd(vdda), .y(net4), 
    .vss(vss), .tiehi(tiehi), .b(net2), .a(sel_cala));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT0 ( .out(net036), .en(en_a), .enb(enb_a), 
    .vss(vss), .in(clka0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT5 ( .out(net035), .en(en_a), .enb(enb_a), 
    .vss(vss), .in(clka180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT4 ( .out(net035), .en(en_b), .enb(enb_b), 
    .vss(vss), .in(clkb180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT3 ( .out(net036), .en(en_b), .enb(enb_b), 
    .vss(vss), .in(clkb0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LA0 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdda), .rstb(en), .d(net09), .clkb(clkb180), .clk(clkb0), 
    .q(en_b));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LA00 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdda), .rstb(en), .d(net038), .clkb(clka180), .clk(clka0), 
    .q(en_a));

wphy_lp4x5_cmn_clks_svt_PU_D1_GL16_RVT PU0 ( .vdd(vdda), .en(pu_en), .y(net036));

wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT NOR0 ( .tielo(tielo), .tiehi(tiehi), .y(sel_clkb), 
    .vss(vss), .vdd(vdda), .b(enb), .a(clk_selb));

wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT NOR1 ( .tielo(tielo), .tiehi(tiehi), .y(sel_cala), 
    .vss(vss), .vdd(vdda), .b(enb), .a(sel_clkb));

wphy_lp4x5_cmn_clks_svt_PD_D1_GL16_RVT PD0 ( .vss(vss), .enb(pd_enb), .y(net035));

wphy_lp4x5_cmn_clks_svt_TIELO_D2_GL16_RVT I3 ( .tielo(tielo), .vss(vss), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV5 ( .in(enb_b), .vss(vss), .out(clkb_sel), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV4 ( .in(enb_a), .vss(vss), .out(clka_sel), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2 ( .in(enb), .vss(vss), .out(en), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV19 ( .in(pu_en), .vss(vss), .out(pd_enb), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1 ( .in(clk_sel), .vss(vss), .out(clk_selb), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV16 ( .in(en_b), .vss(vss), .out(enb_b), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV15_1 ( .in(net050), .vss(vss), .out(clkb180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV15_0 ( .in(net050), .vss(vss), .out(clkb180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV14_1 ( .in(net034), .vss(vss), .out(clkb0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV14_0 ( .in(net034), .vss(vss), .out(clkb0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV13 ( .in(i_clkb0), .vss(vss), .out(net034), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV12 ( .in(i_clkb180), .vss(vss), .out(net050), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV11_1 ( .in(net049), .vss(vss), .out(clka180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV11_0 ( .in(net049), .vss(vss), .out(clka180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV8 ( .in(i_clka0), .vss(vss), .out(net019), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT I1 ( .in(net5), .vss(vss), .out(net038), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(net2), .vss(vss), .out(net09), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV3 ( .in(en_a), .vss(vss), .out(enb_a), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV7 ( .in(net035), .vss(vss), .out(o_clk180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV6 ( .in(net036), .vss(vss), .out(o_clk0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV20 ( .in(ena), .vss(vss), .out(enb), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV9_1 ( .in(net019), .vss(vss), .out(clka0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV9_0 ( .in(net019), .vss(vss), .out(clka0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV10 ( .in(i_clka180), .vss(vss), .out(net049), 
    .vdd(vdda));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_clks_svt,
//View - schematic
// LAST TIME SAVED: Dec  2 23:56:04 2020
// NETLIST TIME: Dec  7 22:24:41 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_lp4x5_cmn_clks_svt (gfcm0_clka_sel, gfcm0_clkb_sel, 
    gfcm1_clka_sel, gfcm1_clkb_sel, phy_clk0, phy_clk90, phy_clk180, 
    phy_clk270, pll0_div_clk,   gfcm_clksel, gfcm_ena, 
    phy_clk_ena, pll0_div_clk_byp, pll0_div_clk_ena, pll0_div_clk_rst, 
    vco1_clk0, vco1_clk90, vco1_clk180, vco1_clk270, vco2_clk0, 
    vco2_clk90, vco2_clk180, vco2_clk270
`ifdef WLOGIC_NO_PG 
`else  
 ,vdd_phy  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdd_phy;
assign vdd_phy=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdd_phy;
inout vss;
`endif


output  gfcm0_clka_sel, gfcm0_clkb_sel, gfcm1_clka_sel, gfcm1_clkb_sel, 
    phy_clk0, phy_clk90, phy_clk180, phy_clk270, pll0_div_clk;



input  gfcm_clksel, gfcm_ena, phy_clk_ena, pll0_div_clk_byp, 
    pll0_div_clk_ena, pll0_div_clk_rst, vco1_clk0, vco1_clk90, 
    vco1_clk180, vco1_clk270, vco2_clk0, vco2_clk90, vco2_clk180, 
    vco2_clk270;

`ifdef SYNTHESIS
`else 

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LAT0 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdd_phy), .rstb(rst_n), .d(clk_ena_ff), .clkb(div_clk90), 
    .clk(div_clk270), .q(clk_ena_ff1p5));

wphy_lp4x5_cmn_clks_svt_TIEHI_D2_GL16_RVT I0 ( .tiehi(tiehi), .vss(vss), .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT FF1 ( .tielo(tielo), .tiehi(tiehi), .rst(rst), 
    .vss(vss), .vdd(vdd_phy), .rstb(rst_n), .d(phy_clk_ena), 
    .clkb(div_clk180), .clk(div_clk0), .q(net136));

wphy_lp4x5_cmn_clks_svt_FFRES_DEMET_D1_GL16_RVT FF0 ( .tielo(tielo), .tiehi(tiehi), .rst(rst), 
    .vss(vss), .vdd(vdd_phy), .rstb(rst_n), .d(pll0_div_clk_ena), 
    .clkb(gfm_clk180), .clk(gfm_clk0), .q(div_clk_ena_ff));

wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt CGC2 ( .o_clk(net133), .o_clk_b(net134), 
    .ena(div_clk_ena_ff), .i_clk(gfm_clk0), .i_clk_b(gfm_clk180), 
    .vdd(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt CGC0 ( .o_clk(phy_clk0), .o_clk_b(phy_clk180), 
    .ena(clk_ena_ff), .i_clk(gfm_clk0), .i_clk_b(gfm_clk180), 
    .vdd(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt CGC1 ( .o_clk(phy_clk90), .o_clk_b(phy_clk270), 
    .ena(clk_ena_ff1p5), .i_clk(gfm_clk90), .i_clk_b(gfm_clk270), 
    .vdd(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_clk_div2_4g_core_svt IDIV2 ( .o_clk90(div_clk90), 
    .o_clk270(div_clk270), .o_clk0(div_clk0), .o_clk180(div_clk180), 
    .i_byp(pll0_div_clk_byp), .i_clk0(net133), .i_clk180(net134), 
    .i_rst(rst), .vdda(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt GFCM0 ( .clka_sel(gfcm0_clka_sel), 
    .clkb_sel(gfcm0_clkb_sel), .vdda(vdd_phy), .i_clka0(vco1_clk0), 
    .o_clk0(gfm_clk0), .o_clk180(gfm_clk180), .clk_sel(gfcm_clksel), 
    .i_clka180(vco1_clk180), .i_clkb0(vco2_clk0), 
    .i_clkb180(vco2_clk180), .ena(gfcm_ena), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt GFCM1 ( .clka_sel(gfcm1_clka_sel), 
    .clkb_sel(gfcm1_clkb_sel), .vdda(vdd_phy), .i_clka0(vco1_clk90), 
    .o_clk0(gfm_clk90), .o_clk180(gfm_clk270), .clk_sel(gfcm_clksel), 
    .i_clka180(vco1_clk270), .i_clkb0(vco2_clk90), 
    .i_clkb180(vco2_clk270), .ena(gfcm_ena), .vss(vss));

wphy_lp4x5_cmn_clks_svt_TIELO_D2_GL16_RVT I1 ( .tielo(tielo), .vss(vss), .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV7_1 ( .in(div_clk180), .vss(vss), 
    .out(pll0_div_clk), .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV7_0 ( .in(div_clk180), .vss(vss), 
    .out(pll0_div_clk), .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV3 ( .in(net136), .vss(vss), .out(net135), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV4 ( .in(net135), .vss(vss), .out(clk_ena_ff), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1 ( .in(rst_n), .vss(vss), .out(rst), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(pll0_div_clk_rst), .vss(vss), .out(rst_n), 
    .vdd(vdd_phy));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_lp4x5_sim_lib, Cell -
//wphy_lp4x5_cmn_clks_svt_tb, View - schematic
// LAST TIME SAVED: Dec  7 22:24:21 2020
// NETLIST TIME: Dec  7 22:24:42 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist




module wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT( q, clk, clkb, d, prst, prstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input clk;
  input prst;
  input prstb;
  output q;
  input d;
  input clkb;  
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;

  initial  begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  initial  begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  reg q;

  initial begin
    q = $random;
  end

  always @(posedge clk or posedge prst) begin
   if(prst) begin
       q <= 1'b1;
    end else begin
       q <= d;
    end
  end

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT ( q, clk, clkb, d, set
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PGL
);

  output q;
  input set;
  input d;
  input clk;
  input clkb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ?
                           (set) ?
                                 1'b1
                                 : (clkb) ?
                                          (d===1'bx) ? $random : d
                                          : q
                           : 1'bx;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_LAT_D1_GL16_RVT" "systemVerilog"

`timescale 1ps/1ps
module wphy_lp4x5_cmn_clks_svt_LAT_D1_GL16_RVT( q, clk, clkb, d
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
);
 
  input clk;
  output q;  
  input d;
  input clkb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG


  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;

  assign q = (power_ok) ? 1'bz : 1'bx;
  
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ?
                           (clkb) ?
                                  (d===1'bx) ? $random : d
                                  : q
                           : 1'bx;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_PD_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_cmn_clks_svt_PD_D1_GL16_RVT( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_PU_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_PU_D1_GL16_RVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_clks_svt_TIELO_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_TIELO_D2_GL16_RVT ( tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  output tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tielo = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tielo =  1'b0 ;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT( in, out, en, enb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign out= (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT( q, clk, clkb, d, rst, rstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input clk;
  input rst;
  input rstb;
  output q;
  input d;
  input clkb;  
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  reg q;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;

  initial  begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;
  
  initial  begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  initial begin
    q = $random;
  end

  always @(posedge clk or posedge rst) begin
   if(rst) begin
       q <= 1'b0;
    end else begin
       q <= d;
    end
  end

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_clks_svt_TIEHI_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_TIEHI_D2_GL16_RVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);


  output tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tiehi = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tiehi =  1'b1 ;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "LATRES_D1_GL16_LVT" "systemVerilog"


`timescale 1ps/1ps
module wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT( q, clk, clkb, d, rstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo 
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PGL
);

  input clk;
  output q;
  input d;
  input clkb;
  input rstb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ? 
                           (~rstb) ? 
                                 1'b0 
                                 : (clkb) ? 
                                          (d===1'bx) ? $random : d&rstb
                                          : q 
                           : 1'bx;

endmodule

`endif //SYNTHESIS
